`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Vn4p7RI/5SCaMioAIWfgUtCbIHQXtlu6Sp2eKNEEv3RfzeFJc0QTb+WsNglFJqklR5XEcG7URKuR
Y6Q6rDxnqw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gLrQDcJza0CPOw3dGOVVBv4ycbKsUL93d5UlVsueJ78cUFQScPQXezBF48wCmSdKbTfhHKuFj5sv
TIH1stAMCzrzEnZMQVXbQuP7IePmpI6wpImEa4cmWFvoZXfSV4SfO0FiZ0v2zVLlK0WCj4gei7E8
nzwcWEntAU4jIKjGKdk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dRJKBaIiPLjKSEGNXxXLziUYgnQ5a6es6jEwSkpVdeGwoTg2OozdYAWDv/euGYX00lJxqovfRiwJ
8LtbaWuQvNkaY99cqrvtQML2MQVXunZyjnhn4FFtD3gRecb8ttrXyev23K9Ykab5iIQ2pquZxZej
bnh5aZD4aHv+dBK594imXDrp2HEpHm04V6184FRja33GjwUYfIgreywEyTS9RoHG09dXVPnGj5kq
nYvJF65SR93nYMgVEvqlx5BuP9YgDyt823gBV3gTZMCK8+hu+9aExvr3kA3ixgQT14jFWeScPH2T
/LxKz0+oipsIXCEPxVqm8268EkEuo62KCHg0Ng==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kT75oxxJLu6S1bclyAxgG4Efp+PO4HBvrSMvQXx/bp5QxNQfelaxgw8H2RxijqD/Ehw7DALhNqkN
zrDilo7LeBauCnvTuthW/L5I2u7no7Myd0+rfJCVbZ2+k5yzQNbU6q75xGZQz8aani1BP00Y0tO5
3gFJ+FdF9mXLpwNZjUI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vSf700Ap2YcsNd60HC1STdpmok2+LLPaOgwLUtHHowISzlv2+9Px+imjI4RrTkr16vdPwZL1bO/W
tsaFGliaz/veqtjrLGcTiOy5ArSV6Fm8WykheqklRz1QmYqqi2CPoAi65+SMf+aZv7nlvjku+zAe
E7i0x5BvxjkwIi2FqAjQUInvcjOT8z/EVsUIc+kBtThm6pnCVZYvpWfWCJhBoTASf3mtpyJgSVc1
shsJ0JdV6sra1cIRmDZmRxPlN+jZ69jgVaRlAvsspaT6Kin4PkWSLXN9o7Dp93Copa9ECJO58miH
Tfdo04JEpL1WFuDCsRl9P/gXVN0t/f/Ei22poA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aqjKiE2k/JKOkskRPYpHmSWE6ssZLBNueP3ANQwfJsR4pWZzmb5Bs9eBPRNsTEaZ5v8te4m6OGHo
GP9WvQ6vt2AfbWHDbpnFz0kcH8bSKnDyyvVFlne2Aa+94xAud+2EkV1eenfHZa8xBuAscS6UXoyW
Sx72Z5Rr2LmiKOzs+rqfjdNh2fBXARESY7bIbu0ULUhfd6ixHY/n4Xtzhkcd0GJTDif9G3F0OC0h
FTTfV4SJ1UFnPsVgrwS8EyozAL9y7GUM1yek9cgtnCneZlWNitXUyl98yDxL7iJfpvd8RP9Wbm9p
o/v/38zX9sJkU9uqzHR86/Np+Oa7KB8f6+Xdgg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 333504)
`protect data_block
4iCmc4HE40oQcF8ccMDamFt8CfzgCgTYNm8NZPapeqY6UaCz1w8RHVI+3dMmzPTjAskS2GiP+32g
qrHzbs7xnt5VzlBLnmyrI0ZDbaWXudM+EfvaMijDQSzpEUlbmuW0QwuMq2wyCz58bdQcXTY56cu5
xsIjJqlrdt4JUMIO6zF6ubCeZl3MFCTHAZbystaBSvXoRrKZdYO2pM5TUqK0vTDBi+y4qHF8k+Aq
980ld718AfpRGSo3R4wZWzwH8Npu2lGkn3cTP/TYog28uOHE9GBpZawiszID9QBQkctf9xBC/Kr3
Kr4BEGFUxAM7f4MHXj4RE9AdCrW+dHiTi1kx/IKJpIJofFkiG5yeFj5jlARhvljnKEUPRS+K2w6I
uDfpk1fsJmVq8Cxn364GesvtxeuZHYt3irwsfD1Q1vFFEDy+OD0K/noWhGA1J56yE2ZJEgFnkehf
HXOx43VWsOa5/BM2Qdp4/58cGhb5PCzV8HE+Xr6XEDRHUZhcyoUHQOuWhYCb8k1qCiV5Dlwvmj52
xJD+cv4IgF+c8mzfP+0tUi6MDOo5vBOk2+g4/H96HPrpr8rEc27dV5YLMdX1gtIf5PATP1fwu9N6
KrPSNIDUZRwK7pHQwSohtcGYY08QktoCBmBLbM7aAnlxUGy9fJ2Cu9GHV6TrSwPdDElpkxvlD9tm
g2AxF6awY0OykZ0N+EyhqNVZHT98YfPM53kC3qFtBDZ6OlLgmbzWvrey873t6hbmLYdyWzVvCsMo
eZiZy+8eMrvO+eqk2vsg+hRNuDya+TWD6p7DInPFO1F2VXdEg0kH6NZlC9Iq9CRcOdpUwXu6oxSg
Dh78a06C5PHYtyhxeEErIJag4J6c0NKJPKiGPzWAzL+rnPr8dfyGORACIVh0i/uOP19q14ayqdTN
aoRAk0hsz1t2tZ7FPL7bXvwxe0DNxIdzeqmyaPsrMgf0YLp3MR/PbgebPAztyitlD0lbyEC/Xf6+
OYMh5tpFaSt+HO4MnK25xrQXcCxyAh8vLZlaCpOo3Q3tuFMo/PDe5dfqJN+p27lsIMfuNReqCFL5
0zabOnwwXL/sdz/A4jXiG932yfzIF6sa4hu3tOj7hatZ+qLxn7JwyJapfxSGNh1GODDEznGw9rHf
7iy3dfZlpfYJKLLnTA4wisyymxnTC2z88yjHDCf8IsFdRXSVX0Q92HiFGk7xqnqs3vjRcwhTYdY6
pcbZdSnqvHxP1UFGt37H4Y/AfcidnujEP1ZMQh7tFrCUkkJG/jTK0e1yCko14V8cKvIIJpz4UefO
wV+YmEHxBMuP8XF8dTIbgcBKg+l3z48DyGSlY0h67rq3FwciODwVqg/Jnw/XN3G7GGgq6Q5gjVzo
Nabz53wqCyAI8NifwHBOP9ixjrHD7fNssC6w53krOHWDETWjZuRuEh8VGUolwdNV3UBKPSmew8St
XNNkqbA0BZYBMSE3p7Q2yNcRDmZuOXgup+87nbljw9ZHhQOSUvm9QfwGSOCiqq4n5eC0sVTGyeIg
QDvY5h/rYKiwJHjw0bNKR8gkLhEOqL33vUHRRN13t+9acIZjKbapF0G7xGg0NhRAI/lHu+gKVHtX
vyZErAwqknw6irg7ge/WXa/xWIUBLSItwv0CKbfStbYcpPPCHpfB3lT/EtqPyewDzqynUWj7jvaK
qkAYXaeg2MogMO3tpNCxX5YkW3H3vUho1fLstRtS+cnyEwBraOUj11pLNnLcIDJNQ0npqQtV7log
7xSyS8h6LS24O/S0b3/Rv5LZt1LQMGu5snY51ukKE8ECGkoJjg/a6uoCS0bu2FgWMWCAvshDmCs5
PDV+/vnLiPCliqDF8UuFTfQLNDmShrrfcCSPRz/ZMpMQ/kn4fqXXVYaRgbEy7vrPxSQMOk7CR1A2
zXtT8yaoM4NS+v6aV4FvyzX4IswRu6x58flKXDbzfYQrF4mphOuO5nW8ycGByBSh0xWu3lKjlCPN
rGHnnFzc2lT++/HW0KS7xxwAm6/r1EUhSpN5u8teICIfLvMumBfzAX3DWvwhuRrKCgYX6tzvsgo+
TCC8mW+gXlP1Q7C3uzc+HMfFuX9sw9Widn05Eet4BlMLJjaT5RGSVIKaTX52BV8/PFjk7pWs43RM
mCuUE/jpXdivVVz434ZvLRBz6j73uSFEz1KenRYDSY1uiNmEI2A5tF8JGeW8IipxKLTblIc6e6uS
ev4nHrT7PbqZiGsoTFFcG39M1gCb2FEEQJGV/17E+rGaTRX6t7tPuYjMgDH+uF9/Q1DUhZv9Ul6I
JrVUQauvBvMRepbyVljrNeQKFJXq6TmXmR/y0yV6ZMNAjSg9wn6aiLXK8fhjQFwEVUasI/dnMPWa
A2tf9chSNXCSM3t7BK2K6PIpQFFaxAUTpfMqaxsAKhjcasorxBsptd9F0exFi1p6lJtzfo5cBunD
Amo4dRZtvHeJqEDX8LVfY7eUnIUAWr6s0MTQLneMwSZ5ZUcCk/tAtuxEn8xDMtYf9XHTpDRSHAoQ
znUuAVXRU+jagh81W8J2KQnLwWWCXdq1EFZO0yptqsa5urCkKP7/b83kS+F0u5rZsr/GBKzpd53j
AtRzlbfXGbdDTlCOZ0QmV1NvBlHsov7SjoE2CK9ksiOFM7ka1RkmV7lcCCNO23DcCSJVsbuvbuK6
0lKXDnGJbezc+306S7F9uU99fALBbIoMzv1qtRyE2VhbPp7IKncYMEWu1HSaf+aV8CbotTOGkctv
TBuxqfwgTgi75bbTKv1Lc8L91oT9e+zj7zi/yZWPRHyBzLIjJMiLof+4HncURCMCJshgElGmDQKk
GyuXFsmNDYpOs6AjvTFCMpwtzdkWXAATk5Huf3mKl7bxmGvDL5SUxViISXaV4eRRY7m69gf/LgpS
FR/LwBIcMh8G3gA+nCe+yHL5QluF5u7sZqO33xoMgysRBcYjL8lO0Ghd+46kow1AYZX9Q2oxO1Wi
/SJevdVHOkKjn98BAfaP9KB82rlKUOIymn7kUFEufaPToq55ydh39Hes7h0h5UZwcvqYym5nvK9f
T+fHOHdU0HclFrYIN3yix5WWFh189bX9P1YfnGWHVxxXg7bVFHnWDKotWjTtUfXvqTBkKEnq6pDL
IBwjsX5rduGl3xJzoA9+6ZtMiNZmM5QptVV1Dcss5pf4YavhiCw9kLxVeNt6653s5+Iv2Ao6pmWw
LAu7EqBjftWU/uzJEuzGvNo40w0BNnQ88eqzoOT6W4zU2A1agjY+H2nGIRW1HqC88MFReaVjXIUo
RBTUuZY23YmYHRFvgdpQJ+OxdTWGFYVoCOSN8KDYRbQ1213ZbzPpNsbdwPGrWx7Lsvntao6dgE9Z
qZRGCorav4AFPY3uoJkdJvG0bE/eKWfB3ByhVw1MthAvFiOyN/oVWkKHO768G8cNoKADLKH1MNiF
Z+XHUioWxvrWSuWFB7ce1v2GChUgPbYPuU4hgFzt2pfLeyQG/TinXyRLItuLqODIgDJp3iMAE0Aq
Px2/ie/9Tt/p52HaDEqWBwQ2PDi58u51Ai9Kq6GYEeWyF/eyyKWEN3/X/VhyDnhOzwMbnvSkkZhP
ri/WUpSgFXW89TgyuY0aWq5WVHiciXep0fOxDoM+VHMTAxET0N36h/3oHr/1AIWO06riVVTxH4YQ
JyOAe3eCS5DvheuHejk0KH3P7wPgIrorIUd+1LuFX25dUon8Y2zzg2/M6OZKGIsaWOadEowI+f7E
y1nKuVMA9VVyFfZ2EdpBL9y1fJi59c1gMYxG/x4Ss+QTarY1uRFBOt9Htzski816buVk5TMjKcps
rh/6dUYWQCcdtrK3Zv7B3mPvN/e0wKScREGzdwB1V+3qatfEDc542stU8C4BXpUhSSv6bxrrWQs3
pufRaTVWVl+PL6hcBcf5cXKy8GuHVXXzxTEd6EDQVfbLuXoJCYvhxM60Zf6lpqVF9pHdqiYMLrax
2TGxxVcmZSD0sGQtTSmNw6v7K6zSV3YyXfdMFa0joC/+J7uUxT2cTbhv37iGEjNlJjdWQIV88xK3
xEfiBf0vtjhQW+MiNVbIw1peW24pZfUT1BRnNg8mWzxJ/KKg9dlP4gkkp0DU7tkdnboAz6dYY87I
W99Orqukh+mSWgGgbFw9JcI0DZHAt0J/uzvFYeVdNgV9v27kVUGWgEDEfKcPhl/RTAIdxKVKUG3/
y7iZhhIyYt7xJZkv5iaHVwQfcDtEjGPxn2wTCEz3tP0e5THtqa1GsT5RxqhlBOrpvSXXuNHEmlwZ
gEiaq9cKSw582ZSWRkdsljG0LAeNhm5K3nmfhDfDgN4kc8FvlWd/Nlm38f2ZrAa1TKTahcNjnXcc
CDYMoWxIHvC1/IGVAkIiE7WYeuqysluckig8ezcLaPiAvRlG535XtHUmQzNDg5iubD7UK7Rk8o7n
MEVa6DeJ7UQkrwzGSo3jryUt/3HTu8wj5iamEVlOv5t5TCD7bVSmLzswgntQNXmiee+q+W7Gzh4S
Tywob/faVZkvm+2Kh4DO2YlFN0ZuGv+GKDC8YbxK0+lb7nRhf2snIVyG3XWfiyQiMfUb8BXpe1/T
StHsigs1S4IkzagDJfX7Bp/FGC7ozCy0Dqa7GXYnB1ozc39Fvxj+QDte4wV2fU8/mXbkQ0g5Gye6
drNKoT32Hmgye0NlkSOMzXGHa+kjjr0GUp2zXEzyaXaBN0BFZqOt+0AmWhfARR6J2O4Dck6nwprn
Ob9nkYiKLbyUfv8f0wF93EkDPu9YmPUgOi/Gg0LBFYLPlB+amH8oGu3hzq30L0tUkTPtFp4ILUkI
GzqPh020ytwK8TqgXUPvJry5BQDn0i9HeiaCnTQJ/kfcV5qpRkzYhEBNVBp+9ze3G3mKR81NgmD4
EYiDhYcFuDeRrT3m3ZrmgqEUKievsFqv76ud56zg5kOBo9eoJhBfowzjSJc2Sm77mx1IYwJPqbSd
5EOh6lW53hsHEZhiiaw0Mq1OAYJINmUIzTHVvaszIH5MlPqyWPOcU8XhhuQzRjC442rpVA5by1c9
GLXF1spQupiN8LoTvcf8hfy6EtK2EfQyzO26SfpMqEb4XgT+c0KwLjhk5G/iXHvXVMufZXcONEKl
ZZMOVJZilkBXpQciTpuRBwoXeU8Ekc/mZCZqGA2KEIZoauxaWGD32kCWGaJY2vFT16d/BRnIXrZx
sfRcZGPcieZgdfb07xNGPDUbE8/FxgkokUckm5jcAef5ePbUUjTRU9mB91KYkwouDWMyDlKXpK6K
mwvqgiZ3DTSCvLw7tNkMRDRl4HoZwX++nm53Rbx3zi42PQEl5A71InEW6iALchsVaXYfp8YqB1kQ
dNWR+owrRygnH2dzM/NNq6jjatdquz/tOQtyr/4shTnZqQ5vN7E4oT1790z+WDQEQmdAhR+KWstZ
Pm9PrHA7lO3uM5iQhP+fDoFCCSdD58xNCMb4hfObmeXntlljPV+t0j5ExmoZUFDcw+8oDs0Vs7ck
UvHa4eVLAi0pZGmQKf+ULUH/fUeGyajjMY6sY0jjGjldWV+mI57tcfVDeyrekOXA7VFSnEUVQLLW
XEADKXK8r8kXz3lKKV9cvwGaX8TC7E+4OxG+/H3bp5lZt0DXeGSZiv6UUcNx/YwKyP3Q8GGNQls8
D36LnQk+CNL6yL1MPgOtvx0Y5N/m0Vz2ATia1HOKXP8lIMrjl9T5iyqbXYzUiGmTMnkjQVRT/eCF
GIdOcaAmkW2NxaX9SFX1HkyxTPCKJabhC/ih4T71NV1rr6Vwa+6mCwN6SKEftVWjYr9JyeQyoUk5
PupsAiSjx4JtgGMF3Aqo5ECFe5I6VGitWPzCpY3mdP+DylkrPlIBFO0zq28xQXldFQb8cq1Dr9xd
Q9uE7yP9mVgwC15Q34/OxQ38eAtKKaFhUdq1chAeMHHT9hAYEJj0IdtplO51eg/TqLEdxE5WOhmc
7DJIj9vtolzA5jLR/V2Ykri61Hic/16LL3rWjLqJ4AZaIBexJwU/gEVJm9Pbi7iJ6Lz+8WYjMIa5
3FcyeQMx6/3PFXC4a4kQYDMl3+b0lNH5PSIXOeW0O3jd6JoX7r4BYB+bgPPxPZ7Dz7d4Md6lwKHW
DVlq9thxmT7KUoUbJFKlMtBFCu2mMr4XILAoRDUXPnFYOpzJG5LmoAaqK0TNhy5SUmhbW4Qh5e9c
gVOWDpLHw4DF4JYlWBdpEEvsH1cbz3MYpmTkrUeKi6PauL97WKhO5QsLkY737N1OUwefnk0PsNpe
4LiMzSMvuJEUVtKaiggDc96u8joQ014aQjvusGUreLsMMPlYhnpKUm+lU66JbptUFXLojbwxOPxl
lm9abuI3jPo92izOD0ysOGbNNeVfecHBooRLNeFS6K49fWfwTZiEJxZcwr+1UbP3Q34H91hg38jD
ZHvXG7TjiA6FIshyWHimZEvBxIuIkLkMKuYoCb5oeu/uCTzM6ZyqbXDam2zSJ/ZPKs4ODNR/v/lQ
SfDwiJnQrnwL76WW4ze5clwJ3Qbf27VrcMeFlMqYomQaeBSNr8HsaiHH63magkcxz4nYRdU7pZuH
0pI+JAJ2pCNGisq6GFatJFtqoqa7cNJbhpwEJjz5LluquO6I8RLh/P+dejglyTaz0uiX5qSzxEwa
vjy61R4aog2vwZQYlkcgSiScQOmFE7NK+7iz+Yn0tHNULKIsUYCkS6Iq9KDwgjBnLzqlYnThzvAI
PrNXXPepZek+y+wFHEh/yJysDzXfraRzjG42x5y2vRHAH5mPq8gX+4vcP+aIAOA7wmrG7jSbhxAo
tchWo5oePrXqRbanGX/aHZS0ldIU+flWTwsgSpS9kqnYlMiakEpU8M4OyCNEnBqsU71kY8nUfBBW
zTVIkAQRDke6Tv9Xqxt4UpBKrAzGrQf3Rv8Mcjzq6Y3RVCS1N1n8dbr4Sgj6zpNVBEuAk0qo+beM
QwJNOaxTLESd97gMtbrrRl2vIjfx5Ir2kgcfA1eA7TKsb14VIEXlAc1iM1BD3svIHYxw8l0HqJ8z
qnnIMtAw61xA9w0B8hIaeNY5UQnnlkpuWFtYI/InF3hdaw+Y7c94cFSUirYSOqZgL/OJXnjPIdX1
GNusltryhjPUtHvg4F+y8m+pihAn8BSjGW/68mi2IXhTnnjcDXzZCGRYFeeqIAJorSnqmmtr3YYF
iIA68iUyr1vusaMKDmNnG25FvjXR5Zcc75DIEjLwTSmB/xK1QMJtKOW1Cb340aJIkLVTUSYy9lhD
TJdAAWok1tDXDrE+fqUgvFCm5edWSUbUkHjDo/dbSF3NvXocnGiIPDm5rMnvABGTssjUyj9oXrOp
WJDXgNR3+/IF6yHV+k1pb2uyAzZkzUE9D5B8a9vrTHsBFPLHOc9XZ4nhwYvQ7e9WYjOhnmJuZzl1
FzBd6kzqMOZFxPpejMuu5E1Njb7bySOz+QYPkp+kH0RXXpfV6gkvHG8dAOmESaRG5STfdkHqTzq3
GhfjdfO1GHto8Cm2ohkWV6Zr5ctUftxgwiqELTeOWnW/vexLRlUcOlpNv9xAWZJ8d+rZGmLbwCX0
LPc32VwoTtNBS8mvFcyZli99tRp+V1de9yszTyeLtQgmY1ph5M2jRqUSz+3Nmb25hEWkSRAgUib4
qIgHuLTZerZbTPeLzoCsEF4miHeAZCe/MKr52kZDSRltakecbcwpK+7sgLXVhlYqR+Xn1vgFaf+9
ST+NeOJcHBanLA2AmJj4/M87tjmPtU+CoDzF19F1sAoRrOSaZ5ejdq+LE2J5wi1UePiB04b7uMne
VS6Zt5Vt4xDt30n0qIqp0heb/D3kR2Cbf/qhnXLKVe7yO0vcjzY4r88yhZW26cxs1jzOWcv3wsVp
Goq+ute0QV/briqznFLiZjWnssav0uH5hcfCOFB6AdYM+cQpARYetq4ldcjsT/+/+ODTObOV75k3
I0AHaQ9mp7n0JxQEYvgb4vhe/9/+/5uruyJPbfRdJSjod2UnOle+4uY3N/lol3t56ugC7UF8HfXZ
4CR1vqRmPPjLkde68LWscpprMaNQaRmGpKfN7K3JC2lS739Vp+g1QAytJ6NQtLaTdYpAID8FoBuX
/d9+oEYUrkA4hQkQlX3olYS0kUXqrMkTevd8RWzEp2euE3mLcKNtVp6/rQ7PBkWqSpNCYqc2KBp3
R/fqGJFF9EhHc0sa3i5Of03kpwWxbHYTWoIxrfVBIXcs5uKqVM72OOmZvysJsbIBdX7S6VtyqLrR
UH2o6AiRPAeHLba3h1zGlBi6Uxa0wcwK75yxnai2tNNPERqq4BIA6KQyBcn526ztQ8TmMA3cA2bU
fFpEZ0Uh797u4Jzgak8Hw5SFfzpTG3WKdfbAPl0wc+L3S8bEGRSNDL9XsVPxd97+6QKb85fdgBYm
H1MqMW2lzRPHTP0NbodBNmukvN7ImFOlwhfz0iYTMBNkRj7rRJaYXgeBRFxdwXQqLnDql699nYHe
uZOZnqwyFxEn4sNw+RnBu2tt/elZrTZNk/9Co5x9e9bA6CNgZ6gUdcKxfTb7PmThhTcm/BHTWTRL
v7xC7b0BVMcyZM1AeTNY8ceIIN4MdOnCnDxbV0Bvpg5n1WUITdAfmE2L3fEeHX2eoQPq7sSZDBci
4dKP2lO7cGTjA3KGiduWPivb6aE+8uP6kBVD7IbgkD7QPPaCjGnCQHmRxAcFXZD3BLAyLxNnwn24
bTr31UJlmsn7aHqPJu9PeR6jJ7jyvRXrGUbCWFp3o9koi8R3atmtKYrsvV/mlDhpgOwWhx9Yspu3
E0ESaLN/NTTO2HyIXTeOCqQHntUC4OcyJmqhRLTQhR20PVaCv/T4iXE7xuX34WIZA7Cl52EERX3S
19RsHjFjXmP0OuzwIqY2lHe2CqpXW+g8v6pyCzMYSuQQ7qH9czDrQUujRWoTaCivsastAhivu3KN
dIdYHomOaKyMHG1vvu2jDB1IyEVEXych9DMW9O7iNNxLM9kE1IpPu5z2d1tbBvPsW+xWgaBep+wE
Nd5jwuyPP0QfNznfMi1SbuUwCaIktWZPQY4+KlAMiQCkBUfi/SeSzdQ6jlDiEcXklWNo+oce5VMs
SXWuu+1XMJhukTPPj7IKH22V2bf6SIgz3vtp6dJblFKPgXJfFB9+JQ+VJzbydGJ/+3gfO+TKuB83
BWHckm4X4mJXSdsVVFbzliiIgdQDX2PdCgYvs9o3/YIJZgVoMxVDrXT6cC/MPesfgePjkW5CCQcB
aZaL98qOn6d6SiO2yPy4NH4ZhESReTKKzmdfDd8k1uEPXsDuLiYo2hc+TVlSGNx/gSAe5pYFqbif
vcvTslArcm2JquErwOSrKMeMvIogTh5Hupigm3E9l02/AD2Fjsp0i+XHNRLMEaJpUPg34uq4gKWk
1KO0m7V4E1fvjzK/lxR4shA8IudkIUYhcjVUNdRxCVIEbBs++lakB2dUWwsOKPJSBuESLTipuxME
bkVdmJs8w9MOXPgY//aWY4Howu2t/j+WRJ2QwIq24VKC36ndqF68fG3bqcUR8LzwvEhF0ljnuL3P
1S5dSbkHiFDIuhKd5LosLsx1nOocB0/71dI/CKz7KKcr7+ZCdJRjSSQZAlMSri0x2DUr+AuHIOJA
iGoT+KIWTcK7Mx3pgvzCK6+qOcMPuxQrzRuxjZ3U0CWxAHMZSBvbBBNwLP+Xr7DbID7HlTf9alOq
vY/pCkMuNNX6OyVsew9q720hzNlSzioDsFDZ9iqCynnm8JDW2RIxMVwJeBKtM2NESPGNfhQmOlXS
lw6OaPg7lKFl2iQ2ujc2fkJvuYAaQfFDZsPohTnIPOHQPkavG2ckI5AKnrsSDQA1OoRIGbztN77r
L7heZaVlgHsRRGOq+NhTLba+BzeA4rVhmzWFr74WOhhGYmtvJkt9Qr1y24Wi8fBVEXgN+6UtuWJk
8Dz8SNZcE8wqitksfaHUcU53Ypv+iXaRY6KlOuYdBh8o9Ch/6m+f+f1LSlefqOjK1Q7BAyDHAgfx
aeVQ4MkH2Fhh1LbGYdLsP1S7CRwRTeJANDMmSPKqFr7po7jABBoha+V/JwfXlDcD+KcISacbCgNj
jRZKbOIzJw4kfFuKJj9KGVpWvMyYfZ8CqrimW/fFcRxKmgt7/tzz2QBQymiNEQG0UaH9zrIIQMx4
/vzBjSkXtFXphuf9K9WPKjRmByQWELo3cRtsq8UsEcMFG3luz8roEC5nfum0eOd0xkR4mJDcL03Z
6sWuXKF4p1kMjcDCHKvjvLPJugMYdMhH016ybahdPFH5jgJGVZUx3ya/hQdFdS5hOj9bX11Vk37o
Os7jOTxZtpvU1MyyuBvZihE4W+eiPVnc2UqGrcuOyx0iZ7K/VhpZzKX2h4qH4X0KE3Gt2ozv8MDC
GkfLT8rQ9Y5LmZdL5Rt8a0tBXYy4ZdBig3EeJO3Br+X35DFf68WdkgWX9vg9cfnlYugWQiCi0OJt
6RzfNSw9TqI4TR1fWVCYugVZsHW0lsYrEu0qnOxGbyq6r0ShRMLu6HwAT93r3DfTBkMOgp/FbFrA
PqjIJBSKxc45uzn3mKjork+/ffo8Fn0qffrCBDWrRhY7dyfxPbeEp8IAEzzSlstY2jKxh0tBvV32
adXiPdq3WvJRxAFEXOV7x6MkQS0DYW5JvArH+HIXBDsbUHahRhKkqaIERGyvdRe2VN/2DFHdcW5L
w+qofJ8kwjzGosLLxxmABs+1+ENFBRpXzebesJ5uls4BHlpsdrRKjZ4dsH7n97IQ114YpXQJuJSj
mWEIxl8s8QF7Stv7v1Lr6prqKD+roYPcPzkw+tYwFQBzNhZocl6Xusv5eTGH40T7zqa/aB4sBQ8+
7Z87wOqZ8QvNWL17gu95ukVTCaj821UQwjAVZe+lShID8SsNRIXDTT4eHXm32WRLv/1cQDrcN3vK
ODnxkKcyc4BzWAMQD8bIjN8IZHqSL1qpYjMYQxaaeSFMqTU3GDRg74sweFnHjEr8U9s5q3k6p7UR
nVOVBfm2WvVUHu4eWrjUzj3ZihpGKV0tVnWnt0rNBNfGDq7OOkeqaIMAyU1FON8kWrpdIwgk6E3j
W+TYDGObihz6UFFJVM/ZksQQZxfOYw40MXWaSs2cXNK3iMCMHYbUcLp+IzIKq/kqVzJWuMHN1qwv
oH1D87PLwj3CBJHj5PaojWIJXr2logT++UWqqTaCR4B5Xei3QwmuA/VkG87xWoWaE7lOM6dBcsHx
PHeaJoQdzkZcs+GGbwVxpOx9zHh7RH+Pypqz/T56T97j+PPZ+9cSJ3ZfzemTRj5QILRUK+vshmH/
ujoSFIxhr87BDA6LEXGJZihaYjZPSKV1b65rhdqdSA302y5uOzKH1RzaIsLeti5iOriL9FKMdNVq
AXAT7d1O5GDI3glUitbdnSpN1vUS/JzXG6LoRNp/VkW2JVPFqLvB+76KIpV4yHHo8Sa+yp7xcsU5
WVoDRwJxBlTEnXJzrWVt1xokUzRpwNMl+LKbASVu9SI2jkWIvGmZas77It5/eH1QAUT+Hugc/qDu
oYxFez78knuQtwcNCUL6ajoSk/YEGK5FQJZBT+CCjE1R6sofposmCeTPSLGOC9EcO0GnmdB2MUYm
4OXCeu6X7JQtbhZOOMehC5/yt7YmFdW0ev/+t8pzqAejhF869zE5tB2s0FFnt77WnNV/tln3SXf7
IyNC09KROMAoVi59Q/udurVbBJOXHvuFPfu1oPrcG+zEOgx0B1yQyJo2eY0lC9hkczZzhJH5wUyd
W6g5zBDHOZ4QuOe6Rj3f6dkiJ758joDZmdwD1dPb1ZicRISlw+GDPzx+0pqhLZ6abTfflZmnxM+J
Duyr/mm4R8ouz0SpUJQgQJDkPYvLYMcn9G4dnZpbCpNXDMKgYo7Rr+vNjf+g3OgsyrqMXcf3Pnuw
9t8KLsax19UX7csvkfXiIDGAe9pPHiw3sYcjwsGxedLK9oUok38Ey00nCDWK6QAkjO+onpE5xaGZ
5VINkBYepmI5mjK2KKUDGgauVwmMXzKVlLfyjWyuBrnx1kgLqhVsjGAIqLCGHSS/Olper4xI/3Yp
IabeJw2MlJDrMCtpvcnsf/rnk2yE0gsVhHpLOWO5rc3Kd0BT9NdeeaAKW1Eq5AL1paWWexcP1cXk
cWLcme8trVrtO4pupyH5un1Wr4ylbYvkbdrt+WgT06wUh1Fs6M8Sy+sDQGlheDxe/EryGu/Qejtm
kMZ60Y78Gn9di7SdhZED/voOaw/E7MpMETSQCuka6jSkRG434w5cGs6iBef0LpR0HUm3zti6AftY
azxHfPYZZqdrEZwH/B4yaL9180RILTnb7JRo4Kc6caBQimqECDCGoH36WlCMiGbp1+1k837YW7a7
rd7N4lGz2eihXDb+hdQ+tWUOu0wrGKRdqb3OFS61+97ribw0MO1F5QEE0tF1r2D+ASB3ojFRXXmP
JElHFj3xmMxCBsYn8QZL6+huZKNnr+49Ef/gL0FeJ8T8XAARIReih06hH81Zng+TBvk+e6JN/4ZT
iLeOW/5IN/g/hDPbZx7Chnh0HeH/mWMGV0mOTcAkW/B7uIl4kO8Em7Sm5Td6zssUMU1bjRU8oGWD
uoouWpL1mrmQxijJEFkII824YcyK/9JiEL7FxJJ2lXMcVNhygWzjJpla+CIUduadhKZPDj9stUYz
N82bRSgE+RHIHapyJUQoahv7RvvMG5MQTMBhsZ7uN1tfjbz0nlmfxSt0Zjg8E1aMdhM+uq2tJELr
LBfxqKwJoGUyZfHngMoXeNr8/ZTHo/jg0flB2QGnFfBdcveLjmssXPgzoyn7BbAqEyQITCbl5cnO
aE3f2YhCDhENEpF3MVw99qvUjq0Tn+QqqJAuZYz9agqaz2f74eUkp5hPXtH62jqoU7CFC3egt563
E19jnFRjtqKCJ1bHMht2JV99j5sv9ddMSKnnFFyiYGt4cIGUIgVjJ5pHqsBz8SmQMSZOmsBlVVoc
Ee8DqZ1RHzJEEH9QaecO+pZjR7aI3Dm54cNwsTgPfQ2Dz5QdzGw/7/4rkrvyvBqA1WR4FnRD9ubY
4sfPtMyQnw5cUDAncRuoN203Nq/UG0/QTSl51swjx8wwREhrHCjg1+8FGIAu8tkcga8ExX50qPJC
nhW7kl5jJA3owkKilFrrv6mpxtEgIyXZmVdQIGPzPHb4snhJ4QcQhxWIhcohSqMwG74qYMAUeGXc
Zc86PQNzzd4+063Mz8d3PQOdgt3XkLIPqnXRk0HrXEAgTf7h7/2dVfsA5KFkaMEI8NGX1QFLDj+b
3IC17szZK6lrNDZDNPIUI6zW7Ufx8OQYQNK7J7AnzkdLiLFr30tKqteukSMhACBqob36kHDpOvOC
n7AUJ8O7RLcs4nuXLqGEdcUYlq4VtM6vOYLvKUlIZBu82bcaJRj5D2ZxJJya6fktyg+xCtUDZ1wD
u7PB1aHVGc1zptQ5FAulGKIhhFzGxugKWXE21s35W2pHvMsPTK4NRGQ/keiXLm0PHqWr0Zf9pmrc
KOGa9tRAGWw8oeTW1b1F4pfRjEGe8lm0QT+TEJ+T1U///p1RvB/G+KI6K5sENSjCWcaqFSNyahKV
hTF8YJJ62lsW5oNeUaDmS2k1RqbR6PExrqgCzrSpHBhvRGCzzZJQZ/UiV1bKsSBxGRGnIP0plPnk
XQNGHAE+FwVbIZxzzcE+nNLNWTSMCC1lJnzSilH/QZK/jGXvaiA5HQSTBlAYcFrNrhbjqQHmCTPp
kocNGhg6J/P3pxWbqvu4GDTcDA4rHu7yWo1Ylo/DoFSSbrNV4tnsJiDuzMwNbIUqDWOEKZJ4ZhmW
xg+VcWHDm3o4l3rOBj/3er1GC7wxirOZDGXdoyjszMziptP44tzAZFOJA/XmOWBEHEIz7dKlRhw0
BXHc8TVozMzchEBTWOkmdTC2zF1qLdzi/CLvgSjIqJaaVdgDeWqB/nfpw0+1KTBZcH6HZqVm4C0O
/hJ4f3Pi4Ic5en8gHrG/O+BcB4Nl0lumywqqbkcufDSRJQLgTVqZt5mPqK+njzJ4YqfalJAVzv0P
yczbGeXKSYHBIAzuPWuOv60idQXY6JN2FnllVYtTYIGHvconkf5JEXHgeyZUhnDcCS3LGZo4R+3G
mHUt/C1hF7y4p1iene+9XJif2V9IWpSIa6TnghR5omyxp3bo2pfT1BcFQf4FLApNctqD08A5jC97
NKFvqvZRSA0nWyC0aufMryG1hP1WkIlEL1s0wz5IdMqXdT9x1Na+hvjXM/wqduk9F6zX2+WhHUeB
wmZAMQtC4nHo1llbej0NVwCdNk/0sMaSbQNQpcEM1A+NdJwA9WPKTfbe3uGhMJHYru2LauXCNfHN
ZmPHNwsGKKs+tRbm1SPo3fuiEgAhU0OlZLntA+o7oAkcuch3iZH0jVlpIkHD6gcFV+86nwHRXis/
yP2VkGd1X5CyVAuXNkUmJMbKl8fV1f2PqGHsmejfhIsCZYH+hu1POiR3k2kAiaXZntGjwCn29SW2
xq+qg7L8xL6HrZ/VL8w0ObhUzpks4dD5TMcKQxKBcyyILFeibnvoTfgMuS/77Twl4PLexvH347+M
glmqiI050sYu4I0pCMQKIkBsaEagzigkkvAUesQtzts6aBTS1VWmK/PxVyiSiRa+wSE17Fg5x8ML
zP7zNsWVTUg2fKkkDobkIxOPdDUq7sDj3zL64X4dudR+xxqv9IF5wwseuZtk5cTVT9KiTDqCUKf0
lbYT4h6FrTdbuXODtUxxV2iOoBMBKvA+GgRXar+jnd4ehsPM6DllMRTETxIpQlqfxBG1kio2KR3a
iTyo/85x+ptFFq1B0i/M16uH2hK9maLkTm7kV1isCW1Bp4DEIwv330HM0JTIwin746ZEx65RmnT8
xq+gtOPXj1NjjbzbXbf/DjjIePwt6mRpd0bmFND8xkd2dS2v+8qWZJvgBX9K5yXs7wRAA8zENkkD
a443JDHqsB++s21kwIzGQoTitTgX+dAvmJe413RGyBhaBdKByjs6n2M5pPEKUoPjgbbi1Lqonc2C
0Y3zO2+GRXrM7qyI4n3WOH51omAjLJbHVaQDPFOH2Z0N7wr9/waIJeEmTMdGzzG+Mx4ieyiD8VXC
acYbfPQvQzlb1R/OVx074J4o73L7BQWmnZKX4MSU12gd7q5uq9iMVLRcJwj11JHToAz2X0bQkoGR
l+QSLUXn2SvQJnKDxX1rMy0I7pI8D4WZLejgua7+MUwUZcfTSqc7MQknbrz2TJKvfyfVcYd14MQR
pqZdDy1GfYij3N2JXP3eITtGXavkNtBmBHxy3sZzp6lImJJ5MzPQwdP2B5uja99cSeSScSFsPzsU
F38cwfa8itvBPdyjpj3f3DaQP6tilj6dbsDVB5yoK0z1oy79/piqpNBGexsSRXgnuIMgqy0+NXGA
QvMMGkJoPCFhravZNPqYrecM8BCjxB4GbsUzqtYXN7t/vVnjMv+z2GBR/LNSOLrYxhYw5gO8FKbs
QOiy2sUKAUaBrZclT+LnBajhpMJFoWrJ8CMrzoOcWnPW11rO76jLP7OUGUAkgISeaRzEm41dPVXJ
sre1oOH9ybIeS7ROjS4lIBIqOQyb1pFhggikQJdspnH24Bv7y/sCRCXQqdSYhNMmr93xg7GBiKMw
WI67Qauc4t02RVLcsr2apg9hOX9rLuudRXQBcNO/HgKva9eUSsyJVxHIZHIEaWkYjvkZGYRnVayN
DNjEYa4yPOhJvEQuJ78DV07vYw+TJ5lDhOAP1VjHZc4kS4rAtHqSojt3XmvA+Ki4fplVhsJPLGy6
hUKHbeU8zUFJeVGn/+fveMFHD0hiO28vGuTtnYsdFqiRDCL2jfMprOu2yP3gKtoAtlQefvNJ6ywJ
05g6i+n46oqw7uVwK1ll8hWQS8Jrwcvg7SBJ6TzgeQdWlMObJOiBE6xdlJ0wvKioM1+fFJQSta5T
msgjbOHvE3NmbjmxHgmSRldvQPYhcJcvw8VGottdSHFCGvf7JlB7Ntv4Ra4AyfSEukiuLdgAZSHq
SZeGPoAgFVmY7O7x/qDTWH9DAS81ljkldxlFH9x7y4SIasm38wuypcfGFpq7uPUQfBQSjz6h5Tx8
gdpaBAtwU4VMNAXNhV7o5coNYdceZmi/p0xYcIp4G0hSRpVWljZzGLbEPBgiL9vptGLXw/inyME4
BhIyNq557Gd631HMg0rRt4d3S1KByvVCxaTqJ9dbdNjGysFx+d+f85QBivAvVaJ2IibQVHloV1Rm
Jy1cfjJXPn7w6G3bVQaJ5Al9CWSmYgOaCspODPDBT4ew2Yvmqxz2j57xwDez5Lx8XsfPOJur/WLi
/bRzWimSTPtIfpcsz9ApSm1Cu7jdpV4fPRaxb2GOBFimS8MLmsWtVGEn8K9Hg2pa/KvigaU2yPAU
aswryXDddBfrQixF0Vj/SrKEC/p2YYRlnG8xafeyJR0OEftZjDiJUyV24RG8zw/TYuxJdq+bXf83
+bpj70/M/UsYAwXCHWMXF/3w52WfPj4s5QiW3ieVi8PlOn5igYF8DSctpGncUS+u/25utIuaIaMn
aknKCAvu4vffPc/J8M/rVZ2qlFldqqNY7qzB44BZpmS6Sb3ShnH/DRXgsAPGdenVYDmBM7DvCBKr
RLHhBemvkjxvkQQ/TpLgxomTJW4mWexilZH3z0PbdichwN7AMJhUclgkII35Sp673i6oRFqfpZcO
YsXuZXtCVRKaWEvthLqtOZy+Ae4uTSzhhMe9h/5KGEABxF/HEumv0R+SiwM1oDx+pWdX0pfGNtF4
pPcc15ZulmHKjdhlbtN9Sfp+wdjeeiaM3jE6VHZCcr5cAr3RMDRBNrGwF2s/9nm/wwSYgTm4T9Or
Z1uxStvh2gmc5BvKCBNgvxDCavZBQn5zbkMtXhsEt65MdyPw2JAE+q2dIHi3QQQ3V46Upn50DjmT
p3fdidAh9UqrHMnI47egQT5CgTcepy/Cp+NlDk3cXB6Lz3CyhAr6roHNw7dETpMEbCnI9Awh/JHJ
lwyXJP97yualF2VrCspLlAXsZ1q5j9/WDz3JCUa7BfBiSCA3+dbpbirCnC7qv2Za3TeJjzi3jy23
pM9b8jNM/tw1X23Vw03YFtpw2X6v4uXl3a8EpT0QA2ZutH6LFHxPYsRtwzApa6T5XXEXQuiirWJa
oVB1Nt52oEzb3l57G6b8uI/Movf2zAnjsbFF+VXj5wXJflhrIi/o3RJVF9+QuofuPTekP06thjah
T1h7zeTvxnW+YM7vQZHwuFQnalFcD6KV0xueFgOergZyZq9EbMgseFh3OdNLiiiHii9VRyI+iaYu
zpV/dICog745tX7+qIIXoxXjkHZssZUwI0iB7mcHHnMX/zNZ/dOA6nQesFBW9hA7Mq8g624UAD0m
Upk8rKXxfQJipES/Mv87WVBIKILiR5ZHgMNOl29EiHNphBV0KRXS2cI1D7ZQmPQiLnZ7qhZl9S/A
adOAd2MhH7ZvJWK2USkkxrlEyRqa6nYumxlRJBo0Feme6Kfo4ae5HOwpNKOuBabvx8HnTsefapo5
c+7FBUuO9ON99NoMGEEbbfR77SqNgSYSRWKz3RuUg39p2aRXqqG0zg9Res4dnkrr97zjdi/NFg/l
g451QlVTIZderzTC7mX+ST4C4UIsu+OwrHxTCjsHFukM8f/M12d+1hIkO4Dj4inSnsot7NrXTmbI
tPQ+GuV7wBNUJU1PW6PlBTrT0MJLR7BMu9xzxQl/nVps6FlDvGGJuvpqYkE9GFBRXUt+XVi7ehsq
ixcjHDh5vPl4T5LpGKOxJCn81xvRpCBUfMlja1mgNd9C7jAgoUFM4UCc191lKDpBOeF3H5dnc/aZ
Wns+W4DCGgv+D6yfW5EcRmc96/+Nj4DGxqkfMmmlO/2IBHPQtmCnUHGqcBfSu27y8KuLoxsWKlOg
xN9J6ht0VZNzjnMx0f3r1QX5tPVDRz7kRtx30st9bHkaUEl+SDxAEZ67mpdhyrEpCMnnDCZ7E9VJ
pmlUOknoVHn8Y1xNqLKDqUUplbRrskKHA6jmOE0Dn3OPY/+l4bvo6WJ/JWOZMwBevPuztwU2pZdE
N7ehwX7h5x0fgMAJSXmU+QYCzzi+oocyTFZ9uBQWRq1V+sfY69piXR2uz8x1YEfp2/GlQgq1Kh5T
t9v0/4aoLk/PAXbHXd7WEEaR36Fo0Ppk499tNAV57VcRMQxzuFealEAHNgpxq9lIP85IXCzwUJtK
JegoQkM8zzoxg30feYbBH3Lc3FIewaXcMHSw0dKFYS1DuZC9KPokRgbvY18mWZNO5EKGxImkzpE2
uz3xxWoG70vinzPftJGp9ts78SwQNfwabERh8YFD3JOK80tPfVHBFYv0nZhleRzUEDNEQ38zIqqT
yQypl5iBR0uX95uZxRb7CZKMpGf3/fAVZxq8vwJprz/AMkWW1SZYjwrSeRcuclwHGk7DSE771ZXx
xjIsingQusEy2EyXoktZMvA9K0wrioSHg4fjM6rzcyzByXGlMtQpZxNsJqLCReaeSjQLk41SHA75
2zLhTfZWaYStqnsZZoGxpC9gMzO2vxWFWrbgkCy6ipPV668CaDGee/WimE8d04sLyws00E58Du1c
CLyjix0BfcIdI89lUdsT030DFjwzy8JWvWbKkz0pF1csl8sQtNN9egub+zCJtqHmTNRbYVwtRMSc
6+JdMVgCxoPo0PddGh/+Ra/SQxr1uQJEBE+xAYmrZ+Q5WgY+oV3DhXKe035uFKlBLtWTRGpvXsis
34FADIOzlrbEvl8EjCC/5V3tEFn4Vwndc6ykuBHFkf44LW5eThwtyqkMvAxWyWqRGiabn3T7XbZu
yHmJSWiSjSH9KJ+v9jBuouotR95EHNo1Bpuo8Klub3J/CxtcM9avCl5MkTCbAV+nW5fRcN3lkXMd
SpBn85M1x0v1nVgAvyaMREQfAk5nxuPabfIsEAWaGStVN0vZ6Sjayy2upowtJF4foGB2KfGCQNN1
3sVafGhM/lc6uO+5yXOYiFacnq652eSWbwkTuOdQ+O+viRdOGUK2rRHkDN1HLTjOChssb6GKT0Tw
A+AmHDw1VoKU6NJz3rashcmJk5LqAeTi9svUUu2cEEcMi6419l1I1Kd8BH/r/mCQzXgnWf/buveO
nuHOZ3IFX/32B4KjIMUu5JFCWjZgEWgSjCW649yaOJBfEgX9JTC71u5+m4wugJmiLPrn0nEa6HbE
33jcUcwObDcaPnTF3CJemk4reKRcB3W+5fBeWCp0mXwc69FLwTqDWk/fxy7CyH4lKhGegwhJSnyu
mgJZG4AvxZJqkTqc3zlgx0WC6bV2a1AQlTFHR8oTHofLdkYKOCMPiggQi9QexoB61qu/j9mbjVbW
BGLwopOCD2JDPw9VeadsmMOCqHblE9XXdPOK1LnEzfN7eocBzFmgxU+NvYOYsMXZ9X7Vm1osCw5k
lfPp1cDLyT+UrUdUoDrMbv/IVSQbQ2XwAzcC68gXDSMuuO8/I7e274YOg/KCwUyEbAlDis0lYZDI
wy9o1BIlJx6CqDKSEytM/pfnvAuy5YMs9LFcnFWTP7Of/5XenkAAUESCKg173zcHOQ7aOBw9siRB
yeFL0StFXHsujlYQDpICDCDUF6eaQLngZcCwpaglTAO9EhGfvZqyovpeA1vN0ntjQqiL64uQARps
Sc59FTdlOOypNJD+DRT6fu37mNI0ITOXa0uvG61hELEVnuWkJvpFGiqLtCiHp/x9ubLI9Y41xb27
GWBHHPbAJUJb8W5wWE8H62qLy4AOC/fPgFQxvtGepp3Jz/n1DL5dY0ZtWv7sgkzcTxNa05kp5VEX
zLBnj8fYQiHPFkAbIn4CXdiM/0DQ26NXwRZzRtcTPHQLGMRx2OLeYHdLLEQrjWcwjyYH1D85PmwS
oyOt3NwyTQ4Zvhdrup+biWEXcKBOKhAoOuwp8+SvY/HBo7x9Rq1gD6GKGAcitzzvYChXN07biqVe
x21zFW58wx4CyztYyiyUGEXr6yxlzT3wTLq6tdo5DYts7W1HOG49lJkv0x5ApZQ3XCN/CLU2hV4J
yrz+lU1BjEqoB+X65SnrOCP8sdD1PMu1YlJWorYKRbnHr8SpFbHdYLzQk9mpS0LGXmHRDR/atMls
gW/dGQD0x3iHnWv51gnqsAu4mTGrWH7oWiydlygs7vr+0o2f77X39Wpc0bc+9qBOhjLAnipaeJik
Z5vmUv4/j1jQjIPTWP52ouxoTwAJXxNoRf5bkTZinrixg9iTWuIVmIzCKBAnSX/sG/B5NlpPMe61
ENYJly6ONoWu7ajfXtaL+zFNMEyXqbJh7LQsb2umhcgHEB+mqW+4y+9VNuIds3rCGd5i9xpt5xrD
VWUu6+oenj0afuplnLCTiHw4LZVTfUDaQMsH6Nykv/i+TKzprJSs1d6byaJ5Vo480MpoZIaZCglm
OCnEgVc9Rl99iEuoX8N6nRtkwmzEO+ETb5JQSgY6h8JJxRfl5x4zGArr2qZU4YjHQhqOFH60sls8
0jDv4lA+e6qvqo7hpEoShn+0tH+MGKprjhoF9qN9NyL8laEVkhR8fzmVTyIyIWF3sBQ0zvWj7/qF
YNagOWkGonF9w/WQK2ppD93SC3oiSaCTAaeJPjoRodB8o0B/RldxaP6aagE2X4mg8mQc49eJZvfr
lqFtBdtn28eycLymh4WE7nNbDBq6Jxri4Meq76EUOOonS+hDctqExpzbNYXvmoqV7ckdHFfw/G2r
6bjTh+kACPGkh6Ubr/a6hE4z1RBLm7iauDr9cuOv1pEvS6Uaw0aVHVyxS12IUAVFXPvYSdUR97dP
3mUuoj8vMK5K5eS83KFOcQeuNCAfGiBK22m4HZwAdkJoK4jxGKw4qJYdOlRT8zNwmSD6PLANHHdr
7Nhmrp3t1BZNJ1WSSrJUZ86MpFZLYpQTtoiunxst1A8dr74sKERw5BdyX+8Ilg/xjpwFqUokJg9O
asOgZO+1w7ujkqnAixnCwQTFKX6ZVR6iCn8s60b85aSp6TjAiFNbCJw7PQjZ7iMv+uIk8tzQoxTU
wWUcJmcWT4B21Htl2Jl+0q6kIIcHyAEBJgJvvV7GWlS0zW7N+tC9v56PqUJLkzpOXSTIBVsce8tp
FqiK7GXyCuf+vmD+OhFYqVfscPDqCR1BfcJOGHYsy4uzLToQOq9UpzIu/3fjj5BfgIPRvGzOFrKg
TSG01w9x99r1IQ9oAM0U/hVKzuMBrWsfVY8uyFJb8KS7aMpJO3ZIGkGXnZ8rp7XihhDWWcRi5LeL
cOQrjnemwyYR7spqN+vzBJ/DUQygF4IsJqCVwl9EmSbTyawc1T9fUTeTuDg6ACFFQ87/RO75UcF+
5WpaC+jaRUHpQlclZlwK7+KwTs9iZAGAmJLiJak68vgsHw81TA2PcZAcP1nZasg+1VT3tcfGwu4a
YdFTayPVOlLI2YTVdKVaBKcxzvNm/BXxU1r61y5aEYKdr52tPJDt3SzxYy+rv3UlnjFaAyL+Ych5
9pCoef9F+dB1UiD0WLh6NUVUcF0+hQY/YUA9HD76YqMIlFStL7z1ySJ6V01vDVHn10bM1F0BC1KC
m3M1QhVAGPyLJV8c9NZryvdAM2b98epbI7A0IIMKkJcmO0nExB9GRx2yegSTt4SDDCKhyFC3Br55
lTjUKn46PRQV0LyAW0rMnVE9Vk5TnMbaekMlE9a5cYpZNY8sPyf1Fn1ubgBgkV7cdnXff/56ERHu
20cD0bvahu1ARP45b+YxYOED7a8js9obs9qGzR6LUiQOw07cuB7mmvSbPv2uyDT0qHZD9E+07Nbt
/6D5+kuOpy5FKW3F2Poe/N/+DgfKtu/kUWIIYmsnkuEwfSlznakBe1kmB1rR63vGHHLHRHkBuSa+
WFLWU+lEmxtkqG2axcWMPMQc0elSHlDEo51eMoUN63o7cC4swyY0SMPSCA+NwAR/dLN88R14aJw2
UUAy5QhMnjg6dEv3uEWVUWSTDrVlzoWOGhsoom5ALpHWU0/UbLuftfAxw4lx1IxBRxsOpaQAa+9W
D6BM1sldFH8hZB8s7nDc3W4pj1/ini1h25vbyGUbVpxT8uHciuzutQfITC7NyMQGpew5ZK5BQON1
rItsGe4XqJaGtmVf/C+yt3iw5XDetnat1oeCUVoNc2uY6yCXVAdBft6LUKkvIj2pwdcd7KVqrjRR
Agqxh9PDI+Rodls4DpWNEWBV5lL9JGqQ1LmG6Sw6J1QevQ/UAlFyh+H7YKHAgmSvskk+8Wz/T78R
jacMCI1bb09Fw2ILGHlbbYsXOCoA11K/lC1Mxb0JatqAvBrW9SwsYYLZQ62o2LKki8aMxikLYge+
wepUiItAUtTGPadSChVp4A2JtY6zUdPrl+s6KYtkpaXYk7biRD3977ypm/GYP1ct7YQLVlhCpfZs
AT/sK1sl3x+9UCj9iJyvWyk2EdJqFlCmIIzM3Bk36EVGZd4scnS61DzDLr+v3k5W2G+YiV+Pekyl
1qaa013FFJyrHSLRPilUzvzjWLl70ptKKrkzL9v8/v4RfMxqsEvEJkSkARG4bREZzuudhT8oDlkY
OxGoLaCnU760gz5f4+8K7g/J4tq/vzob2fZ2VsdOJ6KeF0V4qaPP4q/Lcm6NUgUjo0cgOJmSGs/b
BPVLQVdrMIYNUYFqB+JI5QiPhSww8THh6vJT+Gc1M3eo5t0TqN7AURI+XB293Qod/VRfcDi3cYNw
7zF7dse2Sj8rEJ+FOkjV7oREeFMBr1/nMXa2xHr0B0jiAQStvkifDdGaRNZndG3yNPe9/Spahfrj
DvnBFcEyP9CytSqWBxrSEYjA2zZVcPLWR1ktyOuVwAhQfwJsyTS0BYDiUlMwmO+H42UgMWRbp5Xw
3xSKULbhvBhQFZaAN+frCWOQiNBMPOlKUjLqYh2QchYYQYnPxaCYLBXOg4armQR+KEL7CIy8qs8L
0LFZ3SkJJKgg4DOsMlQO8yp4sMT21AZMPMI5U0uXwzHZLqQY3b09HP6tvU23NaBf2ZnNtzNkCqs4
A+yNMO+eqYBWd6iO0q2YQQiZDq1ev/+hOInoDt5rd8kg1rE0BQ27Wf3stJ1w7fNFloWdFrOZjy4C
HlLPGTrPz//sMZB7eVWCX0LfrlZCJP0bFchXJ6Ky6kSoE/rAqyRaag0aJxFbxunq5yb84bZMIEZS
KD1HrLfRcLCMx1PaQDSvjM5AHcG1Lox5ljcMvTvOP20wzg+gchWlb1y4cI6BK0sAb2U2MwPXTLLt
GaylkRz+pCZhjwfNYeNFXZJFhdAeXmOqMjq0PnxknRRESMqhWQsp/CNghPTb4ul7Ak0KXQYsoVYn
Facvx/Qr+X9U4HWADLtnGwqH84r8cKY68F4mfMDoFzZ7+FLhRgFMINENr34WybKV1zkkJ+NTBjS+
7gj+GLlkpIQ5LMnIddLlhGW12st0RuOoP5+wOggIFi4alIqc/3W8xsAfMmM04mPnhKViKNGBwNjb
VVyzV/fAas8HraDh2U87qgIg3SzXh90/8DW8FZdAnfcosHW9b1bIetllC1oUEMGTeRjz0/+Hu2o5
bvJBp20mw8mnr/vRQWQ9KHM7zJJSla3LL21auiAo9cbl2Wy973vHs/8q/PeyYDaV3Afjaoc0ldTu
aRPJSxfwO5qkBIjyDd6VgSaLc/uMiM7jzEtKfZOzXOo/rQihCPCs+GdQJiFMCUzT5EwLYuyITXWc
YxEGfvybrkZdZMcffsOU94yUAsJNWgoeGn3N4CNaO7O8kjMHX4/9CEm/fYjI+R+UN1bsRVyTFkFr
DprBG15N2Yqk5vv12xNa5CROJIxLJ4D/RFqOt8skWzp9o2HwZ3Mz9Ov+DtU0AH9dVayVCLdpEvhz
d4g5nQPQMjWiZ5CoroTAyNCTaep3XK6qOwtvTFIVv2anxB2/3umvFaru+6gW/3pcyURJILI3JzzX
Mnt1YQaGNFFGw3xEvFuAYLxKv3qGoe/t/99nFJA8zVtNvxVlCJnD+o1uBvG216c6t9AN9WnQ9Rzm
+MaI+Cr/LwaNUvp6DdQ6l7YZLRUBVLMpzOv1d0PrOdwR7eO7aWdxCeE3VJTDczg9PyMYrHUU8n5a
nWYrbG75WLiBLGOH/pq7UrUYQFMIwqFZ8otoDVAdB/7EeUceLnWW+V1PQ47t1mc3OCK84w6WQuDH
I1xWtFbmUehwan3ri9wD6KBbi6eLHDc4hGCpWucrsdjxr+GlBsNJQVEszh4St/Z0lb789aJ9PWQQ
Sz09yZKIRfrBdrmQwrq5rJUWMLtShHGrU+GDrUM78+cFyh4IlebLuMA6RM22sOnO+Cli3zJl5Ubx
0SdKlNJXIGuL9Z5D/orNCwGOWeKEGPAPxPyr7Zy6SaUEUMBk8jwyfiaIdgDBtSd1lm+QBEzdsGQc
Q+LQ2Dd+l61IdyVIXz5jmdhhHXyLWh3BobO2qK2l7q13XB+PY4Lduhux/WC8Y9mRDRP5pjg7D1Me
su0x84bUAMza9PNSdF5ucTibsOr5lrqDn3XpYcOoAPCUNxw5g0Mlvb0YaiqZknK0YsFSHmA/kEOX
dxB6hHRA1HHSSvMSsu14h+PRFhv+CH5SbthmYpmnqm+gTnKxPkfXGNUzMez2yj3uV6Z10rOy3V6g
63KORL3SyBpuAVjv3O/GO8J3L3zhwBcFdvQWhAuu8QXXfnIOoDz0OHi/l8n/u32xyUrmkJKM9iOR
X3G3PIM/BZV5Dn8aotYbRGByW4+VP2R4M+IjPp2P6h4DQbIxIaZI9sElVw2vqcjV6YFwYFb8crve
HQnu5PSX6yZYjaRtkFPXRiFYGdG6JVbmH92AxYjpq/B6Zaxm1KRZ+aKYFMREnqT3EOW/1Ylieu0H
8hCjA1XXmagnKEbs/qZR5RI5+iJD0XlI3MmDIrxnn4181szMRB8QEO51tk5rYFBo5OOR2DOlUXyl
JYGWW7BG4pYWLu0z7AuZBNQInNl8RoImG4OayI94BQw9LsAD2DbWPvsdP9GtEk0ujbw0Jlu9MdUr
RA70f8Vbo1L0Du9a0UBSEdsQt5oDI4t5p+nUBw2BDf3qFYAalbHnlnt9PE3eeWqtjFHFsdnBWVns
osUDk4/AyWfnmOj26NgiEGhGmwVqYBCY9VhFktLTZoJJQ7DeO+qwD57bZnG/a/I8Y3b0k8Nd+aom
M0ii1RrYKtXbcVDmpy+MFxCFGCv1RcZKvxMbWF2f/Kg9gcy37dvL2nRSlhYrHi0kRlRIVf28uTp5
I+N2eeP0WYEo2MWC6f7CO76EJuG+FWtsqf5ybF5LyUnXuXT9xF7dSqDl4gLDIWIV+wmAUn/42rtM
yn9arIFj+0wKELxcFNPii8jd5FwKIELeV6IpmvpGDDyFXy03B1jvnK6piFVRQ3VsExnMHxVc/nyO
DTXSxUwHZAdelUAc0ZgpldNIaJFp/Le2CHb7i9J5O353INM6/L210zny/0jjoen9Z2AcLeDBjPM7
35L5rMWQYo4D9YMQuGvc4ZDq5cMQnkF9dX7tcMkDf37iEuARl03WE0nbKQX6bvv3F6gB9G03GP38
C0hFoamLvBcMa9bA0Bv5HPXeaKapIPV6TmMQ28tDf3OqHZz5TuapaQkRG9xd932H8SEWcIPniqiK
IWFn90oF4IX6v37f2k0JySld3gpK4Sz4MLCCEKI6MjDU8+5vG0uYkDWTf5MExja4sbVgKBkbw8Uk
OoRl5+UMHW7rtx7sYmO06zFUzFsWxj4oz2g/pqpMt8a8q/HHMJ1Ps6nR0deNPffIVPmby7LRCDwP
M0Z3/CmhwiF1KbRPaw8AM1VMqgIkV+53oSEWS1/5xcIsxdeivUdlSO9PRpx4xSgobp9VkGHdhQTf
z+D31tAKVd+KytJXEp4F5mNCqhOKvBzazfneOPka0lb0B9sWsNvyqVWzYxMFMLuV017+MYONt61T
nwI72IOOZaQSSrtV6g4AgVlZdXD1DIQjlf+s+d+OQWlGophJ5mL6i0m0q7Y+CUyjO7Jq0FhiXYzt
f8ue3sX19l2bQkFDqm7SpjpTXeTIS2TM4qyB7GApxc3lyDdKvDjS3e3ydnW1470948LjLnGFPrrg
DwLXmxho5agll+L187nMVc41P86DOCZyrzPr83XsICjLU9IFrGYEiidfqvWCf9biR6nFX39zSI/q
numUx0kLIOvqt67OhyHpVSsxIt6F4iGvB8YfjzX4ToLICskRkB7I15S5nwFQQeO+WsQ0M1rcdFS5
GKb27C/HSdcGOmFWxx7xIaHRjHC0Wf/pelL8rp5tMN6ELs4YSWncVp+4tJkdvT579RpbmFeiXAnD
K3+Xt4wSBAyEKNv5hUMfuq20vWPrl8vqKxLF8AJyuqMGOpB1a3lWHtXGqsIzbYKIpFRbDxdoFNWM
bd1ndmJybWZJAXfZ7/3smuydXkt9BTWFganVhEezJI4NEeBNWT36139esuPvMDPcxEHC5WJgnuo0
gPc6kP71ZyD7aWDzNnPN0ZcyKbd7UK7Rr3CejdQN/uYEmmgDCq27iG4MKKeAdAjGaZDq0qZ5Hb6U
ys0zxJesSWvDhprZXNqlEaT4bv8tGTWdfCHVuw9TmncXmbBTiajizgmVLJ9kyxTCJKOPc+CxrKdH
PboVwxDyIAPlX5DdEygnVTAgT1mqWhBZPUxqSmU4JeMDRAnQ7qWEOqTGp6/KujGXO8Fu0vtgPUr7
QVoRx6/RQQIooJmPcXONixykBVdcZ9a+qbEZgWd5bv23LXp/Q7IPUJrup51r4QA4sRDT5HWSzxiu
DMBnJuK8/jvg1r9sJM5RK4UBNPclkE8V/fHKG3FY+mxMv4QIwAnY/IfH5t7k2uSpDhd1TTUdCml1
e0YnSLMjWysVGH2llYLv4BJVipQND8TZgIbR3GB4jLCGz6siF/+n/HPSmJBcCoqVehDKiAFbRge/
LVBzMpecGu+wOd9tXxVZR+r0ebYm+s+gx/aiy58Wo55jfR9j1oKXhY/Q2pEfapo6jYOKEEvwPUE9
Iz433yMwNycsvkJku+V3p87S5z86SiA2KFH7jARqdb4qpJrwJoyD5JNqaY5iPEI+hGenbnLFlDzC
Sb9X/rYiVLAU4p9nW4EzCFOnzEE9bMuhKY0HYjmyY25kDna2Ru58kB8hGW0ySyp7NJSNPy/NX267
aappKPsBMMgsFRelfWnU5PLZhG+oO2ZJvHnn80VRNaUJm7DByTmY2KNPFozCa0Bmii5JMYnXf89S
8zry4n7BcKKxsAkdKVWXyjKggnLcduBS5HK8F7im29vLglSoeJrfToL3eLrT5MjlrltRofjox9lE
b6tAU4PgzTmW3tOaWUqSRLhOf99NoatTYBZ1zIqMMmX4n1YnK4wsSdjLhM9M7pHol+tPvg24k5sD
Fb+ztaZehg4yNcX3LvgtEmwOgnMoNXD9ZYx7gmYlAKr1X1QMMMRwVjsm3dva+tP97TOBVTZtG4Rj
Ull3XV6fSfNht4mjbgIlFmTPzvm55tIIeq3NlDg7XaR/p/C0O8sL/prqk2eyDlyJu9Xti5Ly+ej1
ElTgQuTMSbV3Pgdz/41HTU+NU5uCl7RQoNpFxiW1mN7JrvWkoRK3d1ktk1+pIokKKYFDoSvkeLrH
36Zg8p2b9CYW9ns/lCYJrT+Ugk82gCmgFmEU8qJzl9TtS9wuh4PNsPyZalNw9hfgwCt6DZQME8l4
zr1iHF5ht2Th76VShqSB9S//OrcYK76ncGeqvUSLg09wOWuw6i87nFZ9NQ/dWLHsZrwK3O1+gzTT
ljV9Z/NF+SKIgOLIaiRR1NBWpqhPUvq8BFiSbxnWjAWaqJwY585EryySYdOqC090+3he6XN+s9Cj
14JfaJpS2+wo3kouprrkoYPuAk/kn8htv102iiDQNqJrM5BKT7//5PV+KsV0miu/mD8cjsiudXMs
hsxQxigOd+KJi/bA1kSpwUf40DuQH90Uu8mCYOYP6q6uifVZiFN5wS9dxv30c3xPEewHD7ZuEFMy
kp5dBZSAdWRx7Lv2DV1FuG2rtnF7sDoswlER+8ffqyBCSEh0dBPqaLCsOVTjpMYER6tcyA27qJte
07TvBmd/jBEJ2fSMBnCQAihLrseE/j+su8KUy3bb0Jp3v1uLWyNMBnru6v5FJc6JrihnFj20AOtP
XXXx1xBwsyzeFWyay4aNZhTTHydRwLyGlcvWRqmTNhZgSSDlYDbw6/0zeHlLwNPQyk9q6kA7QRdL
+eBeYhimxgFE4N1Tyk8tle76CUEDJX4h/W0YbEb7/DOTWvJLOdnkgTDMHCCZB6SctsdA7sWVeU3y
8fE50r5cpLaf54jPSK5zRZRIG6vf7d51F+DOYRUV0UzgOjC8YvUWQ6IZdVdop/PuYvXX8v5tiORz
aQgCjyAFuvMlvcLE3fp//FSWgo7AL8nMS+ESXUippQkgv/WSyiV0g6zGOEOu8L53/lttrJOBA3x4
9AeUhi8wYQNXV4vUktQOPFoSbJgA4FN9EcXggRHG3NvinZ0xmE3GAJTCLwkADknE5LrhCzMU/ynB
3IGwk7UgxVoP3NDDHbU9sMv7eg+AJh8bU6xDhIGfhMmDzEAWxaY1o9wS5fAzxQKi2xcppZJJ/Ivv
mrFbp6a1evfNLqHcopEyWqaT4TmAHswQj7MpPwU3oC3KS3c682R1cbSEWxS9C5UKrININtCxAeI/
4kzsJ+GMEhovSJxqk9qNERMxbfW0lveGodB0xBprc0u0aBQruBz+yJG+KCKQpnMLIhDhkdf8z4B/
1sVewjdhG9tq6X61e220o+ncQmoiqvf8tDY9mM1XCJsTJTwR5wsEyeBSG9iLZiTtRhYwkad9pAMM
dzVGPpMA1xhX8guXq2WKyH06TSB/9OKXNqfIj06c9ehIAmKZGTxUE9EjYwBVXHi9FwvbVqFHSF1i
Z6MT0fv0TQE0KizTLSNKurhIM96CF/Kk/cvP1/RYLZeB6zVE72RuKehwbJ10YA53pvxHMLSxlG71
PDFKcDTUnkWpytUakuy2w2h5xMAVdNU4+IpjIOgnXTEexv0POQF/C1Fe0x252BX40j5BmLM9tv6j
NSEaHwcaIKVLXGVV2cS8Do5uSfBDzkHKxLUHCUiV9nQtL6bMAn4/3FhIgDgJKzI4FWgtKhrKP0Ba
ATozNNzCrQPGe89f08BCUaG0axhLzWj7RYtXlIp+7apMszgU9iBvpXAOnhIRuRbW1fno1jJEj0so
fqW/y6kOFg6DQaQBh1megFm8Ei6RUryqU5cBd5A8JqnGl3YzM83blQ5Poa3f0l8wivBNPAWlMIzr
vsNRpbqWKuE/FutGBoD1px0hSyKssRv9S6buXfFZKgOUxA19u//Q8NKzWbUjXIuQ6yrNE4ioHzES
3CdLSS1Oy9jO7/UTH1+pqdx9iTK+g9oUVHj5CipDwYA/2xslxHvIhFDS1A2eBPbjMl36Lgqv/x47
y+Gj3dHOMQkKDm+I7329b0/mRL0u26gh78tEIq82weARYKDnkT4VbJVvSt42yKUkxGg3vMhCSkzW
ZpxD3iAnLBv4I5TbI8S/sJW8N4o9pAA4bGfkIADf7BdnQquepf0bMn2aeMBWxH3k9UWsMBo+zVYu
i/rWEFH+Gu32VFJxwcQv+6g5FALgX0+hgafRnTsAmg9B3GIXcF5fEKe0X815OASGO1QQEGVmRIVq
VeWUbg4qSIPw8krJDNkZoSz4KyfQvOotqN5A3lk4rtC+lZKXO66B87fOBtH0A6nZtcBca66pC0Sg
/udDkI+ebpouJ8L9JG0eAhRKEMdlJkEMZlHdSqWDpS2svZUoffRi+20pA84qbOZ8JgIFZQwXE3F1
/ZFoRlACSG2o62dZBmkQFGJJKxUR/Qo56S5nbL7mCaE1IySaYEgGK4WlgX7j5kd50IxUxwEcNzYG
a6QC4XKuXCteeAxWbb25I8BaPYms4nYbNGnXQEAx3b6QKJNgsR3ARdeC1CyBsd1PhNjGnzSQcVQu
fbcKoqgJaz98qAGMuuBiDzRBQnLh3xknsHQoBUa2cZrd45RaDAU9AKmkELJS20ypX4C3gMqEm8Sy
Bso63FUKExW8rJlJYULau/C+tssOxso7qeceacxywjgeAie/rcJH0oSb4cdr76f95r0E3nS6wbnf
26uLZa+cQ1b7/J8O+dlFkfL7DVxfoOB/4Yfk7VQ6e+TSzpF3SbFMRR78pbQSJ7fwTKbCNsHxfDTb
FmfAKmo0+96hOpoE8gtJnPluJPz6pkekFpvWmPJfZf426lr6O4vhuowKns4d5NM0mG/4KcdfwLJZ
6FMwlkvLsGXI7xbpLxsPl9Xqzi0+Ert7GzwjGE9IMXpqQiFB09/3oWeon/Wb13D/ve7fBpOyMXfx
J/7HLH1ayOjafbruleLmbWMm5GOjreHam7syXYEzZAA8yaIP//WjujrPNzJ6G1xREo4fcs9Z2NQA
+B6SOVpDVdQJtBkjHQWo9XrdgynvgfVbgUJK7u66iaPeJPUzf9wjed3395BurKznfkXADgsA7qdY
K3V726ep2Zg3onY4fq2EqzD0kJ0+EEusyIqlfGZrsazxKcrswYAaRCp3KzuHGZTC1lV+76eszvAL
o9ozpgSnUz8hipfx4OMQfF54cdCdF7M7brbxGJ6f9My95jx95LtIEAI4YEE6DmziRTaOObW+FJ8m
aNsbEkb2U1CSt0kVZgPn3DnTCUYNiM7judxKXw3YOAw4VOIxh3owi6AfpmJM5rO34xf8yMqQ2cl1
X6AQUY/9to0+YsKKhhoM6ZataG/+gok6s0zE4o7aqlbO3OIo9ns9LlK1uVsQFwZ24JOcDVoTt/7u
bcPX/yvwdIE4N84SDSsApz3UJBmsAasNKDtOjzvbs0wavxZmjUNJlssSWlDsi3Quyl6u6sN1YbIV
pMN/Ge9OcWyGGwKGxF+yXKvLFweXDfZAcaDR+z48nDu0yK+BtHVwNcs3a79nyr2xcSYBRDjjLR/x
TjUHGiKUN8zDMIWRBsezojeWpvqsdI9ZgvOiNq2OGeI3ZuGmEVg0Mb/PgBZKtoQemAY2ZqqQ5fah
7p4ycXlMCvNnbRM/BRU5yJlDhKHx/kVhImn9ks/9fyIOBxPEDAsiIVZeKcndar/hefT8AcNNcaaZ
p3HKvbMtAFquuPuZwkAosqzdeoc08nHfSOtJPP3hIJDINWbCZsH6OoWjFOeFlrg7GowFCGW6P9oF
+W6kGStXXfIB7h0EZHluxC42wbHDSiK0HakcpU9rXHEJfO+PKJSFyy+MrNNZrVmmchaafdJdP2q9
NPD6zpLzx5ZjfEgcs3/ObsgNS4/jnBbvMCKSPit78dTn3zhYVN0ZYucRj2VHycr02rA3OWop+0cR
zUPGgXyeRIosReYMRA/qhytcAwmx83dGyMZj/c3lg0ZG15YjLEL4L15a7l71em2SzMZJP2tRs1Vz
zUe4bR1ul8jRUgUQsP1J9XtKF6aV7A9RLBLvjz3NHuJTJzWl5JKr50bEM/IK3Pw9druO0pNZW9Fl
0kSATWvjxjhDnnmXVqOoJ6XA/dUKmEZVA969O6gkSMDFpUcAw1LOI/qVAZNw3JX1E1EeASxwmiHz
ks5/Pw8cp4XtTacvRqR2DFZVE4XoFjLOtd5PCyuBzClBS/YE5P36+HiWAOLc78nFOZoUCjTJQ9Si
RWbzmS+QmnTDsH9kXap5rWsrFe5kwQdYFfiNm/ypQWRbw4IlgDxyf9aAmalY5CSu3k8uLVJQaoTV
NFW1e2v1SyPrGJoe85E/1ynmjHYrulc13tzjcdLSygm1tkw/veD+mJHUlvpVpKxFhcO/jdDAh18W
oM9HRhHi83MyxDWMgny2RJuwRespbZGJ/5WJ7Pizh/aKSdFlRcyr+K1NOekSZTTjWU9TRQgRCySY
b7FQuTUROtOL1lJYt7dTWif8rRE8KRX/AgBfc4IsvNfdmDjVlX62cjjRVnCcjSrulDAIY/vyy5L2
Sr7K6dBNgk/T7UaT6KPcFB8w7ouNMBRLcfvEwf/igW0d3KsnZxXOvVB6/7cZXryQrcGKujJS9RZK
WkZvlhfCQxw1JiTh3fsI1ClLhp/660YNP8GRYvy8Ljle2phamKfM6K8UXuLswtWEdqCBy1XbMc4b
iHNf25B6LTcY3QOpvPQlzMvj84K8VTdiiyZrPFsPfadZdtyQaJcSDhbZB+tQZEaV7RhJKHpWlvD+
ZYAsSStGy+qpCEsSPsEyCvQvrV0flVgUM5WOCRp0wRlaxA/R6NvScyQPK5A1z8+kmXkCZhRYXggR
Ai9sS3VqDjIjjebeyU0GYyHXrljA3fX9hlA6eIuTKrtBPvRQao3lbYvPxdm3tR08uzpLQCOWob7A
R3myzYeCJ2ZKjqitzErUvDhqJ5W3KJVrX/XYC8rYjvK98pbIrXmEWI9fVQVc92tXYfGEqWxcwARy
kyf8TXzTahbjKgt/HvKnpx6rcn2AbXoeJ3M+25xWTRyEuvT7aVgsFE670hSMralLGT5OPUuqBK0B
DWxeaOPdnJlVRtpkQBYfpZQG4Z5FeZsF1xpU7X3BWX3daP+zoPhqzhghMFn7yk5l4euqH56A48mD
EnaJCCF4rF6/EeIag22URwNq47l37RH3FrmGsGCxWnOvhTBHtQJ+nbndct/uIqGzNDIkqVsjgSSq
ot5qTsSWZMBTOFxZeVn90DIE73aypNEkjHdH+mLXz4+HMCDd9mgS39pzuY0j0G9+GUu+gYV4uLk7
tRKtRQZJ2h4L8rQBmPnEa9J6RB7k+JMYnCv6X1rfq2JG/TqVkjjy3hSjm1ktLZIaSusa+PPje833
ZYTZN9cqDsdoPgn+13K2GhDBYwsylfJ4QtXZiOjl4GXwLssbdQQPU2VG84Ml4dSVoiXGmL4a7oWA
pGBSDPsqH6neLJL/ICTpX4VXIDUBayFe2U+aP+tePq2c54ToUu6//++uw7pnRU+EbS5mqGDD+r2y
8ildNkNUu1axgHMETccpdGx5yIBlfdaRu13yKGsCOlP2Hhbn7y5Drd1xBDL/0VswQ9IXqJy6lHhu
l6abJw3HGsdT7Y4eQ66hx5Fzk2rnWFg+lc7bosRMwOzc/ZtSES43aNRMiLKXUeh2oO2GdXc+VqiH
CEykWU/luvkaCxG/5/upATFK5Swn0vA8hwxOLMngz7VCeVT3vrS+x8XG8Z9u9kbA1JzD4MhrjD5V
Ien+FIJwgUdN3FYSnx+/hNlHub7OQvKgpqDaZyXR8b0ooXT9AZpbEAZGy7BmFw14Az+EA6WdHW1r
bAUP37g5bilLgimvg2yviwjrbdv/Pdmbcj3h4qpuDWfTEcM5KPvAttfMK4S+RZjZalV+9K+mYmrx
qVwGNU7BEvgTHEgTUignxAb6xjYRDc0XKclOEJjN7EbhqhODkE/37e9k8Pf+10Iave9hqoDeyVSW
b5mpvYzKRE3stUrYVY/4jDm8PMutMQfW1Xx272lCWdHOmOV+C55Iq5EWX4uh4+UAwW0a3jSM6TNH
5HPJPoUtp1QrHOaAEzmeKuZ3DxR4h/NHkbed/RDA5PkPrAg8h2Dz5E2QUszcfmLasea9bzhSXHkj
3vUd9i/vxkSi4X4fc51EDZUUwq2K/CAxTGOD3Csl3w+TFvjBTfbkhfk5R5tVCgMfDrNw6Gsvsp1N
iF9uhoQbBUpzDl8gkeTVhEHS4G9R/zr3rVXQJNO/JR0gRomSpGUlQyg6AhoOYhd61JoB/+3+t9b6
EszjFx8O/FAoHzK2Us6OrokeJecx2yd0MKH4q2FZvq75H2uyHGJz5V820OOBqPKgsmOD5io4rPn6
lfflKAZVjoBJ/vub8xC7l9TQsUuR0LFxj3+HpZvhj99KjBthcHf0nW434Qw9YZsX9nYSZlGKJXum
UG66GwlpvixDUamwLSZBejeZiINvKn3uKfzRQHPTguh9koQ2dF6xitpJ83V7uo7oFSTfNcCEdi3u
NARVkT7DsjChuDJSh2A2NaK9N8qe4RnaNd9Ib1z47hkTRBR0KColtb9aADw6DZZpETeMlGUYsKwX
07QBpRE2awipWXuKbNrV2qkUxdfhJUkzdMO9UDca4lAYlCFKALZK7tyLlD3kWJSKhgm8g2Xzg1YG
WUtS/8CfKdhuRsAJUaS+t/ysz7xF912MKX1h3S1RKCAw2Y5ymFIBg5SP1jmH4cJKXEtORBp1rxUv
JtWWNXb7yimUFunY2IQ59lU1TIz/fwfy0QVywf/bW9MgSgj9+cZINVrxaeOY32RBoOIkSBrs4eSI
4zFW6o8Mk2KLAVWLfJ3uwKG9wnsgN4XP1oa3SS4G8IUJipAZqo6Iv+4oT7GLHGErVFMn9jC7ZUwZ
qwjg6t5IM255q9MdARXbBvRdP0+8g6OpV0AnRpBb+AUDoZX+wwTcdL3MRY3QXQLdpPVpxtkIUstv
y+C7FI+irnb3kEjBlGq17VCnhw9425Xymfp7OoFIibxKLDLacx5BdqYZWHuby3AM2RQiMEGpDOZc
S52Y784Y1eOpVhrl2gsChMoG3P+vkKmeaVqzY5p/P5ZUViJWEYvK4qT32Srz8l/FWx8DxISWwwZ2
BctYJmsKLwcjrWZuDvXnEvStpbdS0UAJm1qzjAGrvpA6u4XvdBbJBxtgW/AE9B6k14j8L2cvqJkm
IDJida06cohGefV7YC811JUPYmDcbEYBijW9XxwgC/8gYnPklttAu9pOuVJpXTF8hUEzpvZk1kA0
03lw24FbkcHU9sASy3H2ZQp+MnxjPpZKp1K5q/PCbsHskcjnwIIM3lE6b8FxD+zPltQWa9pxR3He
B9ejNMTuqB7fSttv0MhOMWhkLiVWyw2cy0QYstEcOL7r6I0/6d5Hw7lVGcg++w6Uh1nXjK5NMn2K
WzM3Bn8rqhOgT12Q+mYWZJQNCWmuGoqlkTNkXRI5CvlY+31gD9fgB4450+6MdIQwpUJx3788/vH/
uiYxFSO/XZBpj5JMVYtK21lNp86y/DrvQtwbPn7M+ENJjLxECXJwj37sntgGlsoxmJuI4AF6SBmI
5B19J9lNWyglj8OlXagcWYW6ggxY48HfxXK9yvMSQCwTMK9mGPaKBWJ+EEDw+t5bAQafukhnui9r
Seo1KWYtdM9PgovSPIAfZT9kV8D3J2iNvQ2WPrk+N6KLomsim9Ew/rq5Sn1k65NwZonGqMAY9HP4
+9VXIEC95SgTS0CUoHyBkXD1DPKGuB5ncFluKvkNX/VlLJdDM/EvDDyIMx2cxt7jAuR7K1Xa7ywN
vNzNGGWeGnIIURnAisoswTqkOsEQGTFQyNamUm5y8JR5d1bwbI/OJ+h9Wssk/ekDLNm/GQ+e03Gh
Z2cF7iOS5KtiI06be4F6m159xCVwiFmPgb/PX7JZM1k52D6n9o4jR9Yt6k4LtD1A42wm9jltHad2
aLeafJgOXKcPqisk2rySzhfoQDxN7sYAoQO3CbqMRrtv7jmY3QP1A8jloteCTFKVPRIuQeRLKNng
4eVTLhNl33HVXKXqZhh1T44pOBommVGfjgo6dB9CHWKhI9M5Ed5+49KnPkcdmttoI4yt8opfmmZe
yxRMTDchJdRyQ6XmxpQJ9gVEIOv1dQeMIprbLyMM62T4lif6/tpW8q8ajUmkHxs0HgoIG25ZbsOs
AKNr1hwlkkXASCBhkDFZUoWdizQu9OTZoNevVi9TGB5xjVTwpMqgLCzGAt0h/PuQoUCDnGFmSOTs
hAC8HYHU5bLQ2b8Y3djKV/gWPVyYZSLq+x8fQU5PYKRN8YmVsfS96h9pQIXg76gJSrB7l+N6oLxi
9b4pYIcX8KGk67APCXSOSJg9n0hSQIO1v/9Cm9rSkFbpYpSBf/B8BVHYuDkp/LEOlCq3hS9Dn5vS
O90petUxDb6HsWbmhjiPvgFWYWMc+Z+PmnTPuCp/ns8jj50RML5xUicfp9hzJ2qrEfJLNZ6VX/Ko
BB5OWTRpEpsmcfWMD07J52KKIv5zARRTgtvf/AOTvd/pJJ354vozk/LTfa1B9+IR0q46cHUHthkw
e0DNV+AtUgULx9zJopMfybP8sGVnccf8oFLiIVIwXcBDXfk0EXUt3213R+1sLbLb1sOVdv8/1bSQ
Xzcs9/ksqtZXE1EjBghmAn4tHxYEv0WKLy+A2bmspbCog36vCmbEhW6d2WiaguanZal4j32FICbc
UEEod9pTkvq/WXXbvbEHrMfSibrINkkV9trqWQ8XKog4N9x53TQzYdsKVaWGbvLDVaHhjZMn/uiE
M3rL+Aj4ZzCRpu2f4mVw5n+CUqob6vjZPv6U8xa64tKfn7fTP2p5Swl+tmvxOnXYvREfI8uwsEKD
obUEaHoPADpwkkNutq0Ji2oWxRZNfQvyJEfGC67YDEENxqv0M7KJVKI7dTn6KsqvmTtEk5081/7K
h9EwqyVuvMCcUOdL0qBrY2oye/9QOu7oAUvj3XbGS8mTGjXmNBRxrERckEPdDojZKf2ufwCNTpMV
JySrg244eoiG0izVUOL2kS4B24etYha4sXm/98NY/ZLa2hVEXXbaHEXQI96zdSuUVIWnBfzqI/qU
vDyLPo+NKmBqAkCroYO5O11hjEUVIETmwDs68hThXF/3unoUjtoSNN0wCKHyBohn+abFu87v+bpG
qZlF1kD38XKMR5o8vv7YaDroBJDV1xmrnsN6CiJiHHbWLkUaQJFMm2d/1gXmijSXK3p/wybmKEpF
3rYOHwqklco5Yr1aFcjTn0VbpkgDWaQih/Le7ysvN7Rg8kTfEwxtAnt+Z1OXRI0C74YK5eHhuJ4s
NOuSbYbY/CgwGz9frvdgRDo87w5yGN0pmwe5qzIYAjAb2t4s192rV1sdFce2xfJuM10awzQWaRtA
tqIL/8zyn9MAtfYbb/HRrkNqIy1EL53YS4awFSZ7tD2zyYVl7LBAxfohv1DRKBs5ZRVYOXSKPugg
qEak3jyoEOcme5LBDymY91ZVAY3qfYly/rIH3zADQPcShZGIm7WIPgZE0urJgcvNInx1yE6RXstw
N0mK6nZuetQWRM2wneu2qF9LovpvysVEwzP9J8j1266JsWLIejmInwyhkqNNwJn8IPew2ndKL34p
+BurDSYldkQ0HpFBR+V53mFkp/h1WLOZ5HCiBLqJkgAjseAW/CnRByl+tXLMqp5Jhzc8w1q5D6w6
irXsJn5mrRK4S7HnrzmUML0m7DHix3/MAJsvce1NPus/WKu2pXMZLIc7WKAkYYCtd0pX0b6uouI8
FY+SbB1UCCKv77yRl5xpQ33kcq2po4+H9efcJevuOeJxNBe8yQUtXVxnJdl7fMas+fElRg5mORps
juxX+oQ2lOyFF3Tc9QBQFvYTzfG1uznV/EwATNoJD+xzLzSjxO0rH0hcMi8MtSWtouso12TtTEc3
YeNP2GcSM2N06LQC99IuyeyN2XBObr9uVDH0ZAm7ZKTNVgrMzsV4cCl54Bq5P1xEQFOfT/qC4VWF
zD3X1FGz5nga1Lo28Q0iVKgMCZ24VWUpk60VA2Z798DyS39oSbNNWFZT5LzZH90mXQ9S+ldedMx/
GAtdUJnorMRf7GuxMtq5JP/8rOkZCLjNrKQ0q/Yt9LSFAcm2dd4xAnOpgvMWT4EYDAt990d3NOU/
gP9eEm2HQz9VjzkKvg96m2IQ3wcbZGm4FzwSgBR3JjZDQz+drxMn9s/4z1oNQPI3bDeu6owrtlJZ
HhSuPuQz2Qb+XzL0xT0Lk32hZ2qdlpLzB31fo74C+5tiafYV1MfkEfe6Y+6iG6nyWwnGXDsaVg+D
Jn5SSsiyNOynUP6eoKhG+tyLAz4VjW46GXupf3j4RfH2aErAQjzPFX+XSDE/lKk0JwC5ddlQDzNu
WFxNsKuRrox52velX48FDHypfSfXgzrQnLeOpOgCfzb3tvSGsX3SKPtw+ddDBKB9QdC6jreRLWf6
6h2VDmYBV5dY4Bp3THerAj3SZqJZrWyNH9TaAL0YIBsgryqZVX19E81TIiO9UZMszrtyR1IdMpJm
YPXxJ7K0PdkiplSujt0tBLzM35pfYK1BpYPJJSi59phAnHKjcalo2JEjb5tKU+sZcwr6wZgf3G+K
eXe67zmxOhgDpjm+ZQ0DYcRneWWvfLymqgXhkE9xLu5mU9TgHzNPt/rSEFA0FZokltgCAMgP967y
dFD1qtjtnjOtC1zXOohUR1clYeGsrEBsGspGzue86wB23dSB2Abt3H34MKJdkLNbT7J7MHaYF1ir
P7bFxOVEwl586sTKh36rWJtlDdlfMpQxWEfS0MUV4OVC+y6FG+ilduhZ3A9ctWRhQfN6TvTuDmWy
Gpoy4meGkAfDimJnuIcDX6/gwg7q1+4u3vTTHhqy/oXZV7uMYKrmI6trtOtPxopVH/uF7ZtqJkRV
ClwgDJ0FCpxU1v4CsjRJz9mz946KYAJ6POGrcuAD1mQ51rA1XaRp+0+rsiw2Tlwf4EEPF6tMbwTj
Dk03hZ+rgNAlxZN00EZO/0B6rmbTZAtln0NKnqaJoBljk0qRWeKDM153Afy2AECEDWX9nSh+aStS
B9COiKrelc011Za2H8eMBp6SVl8VlLZyUOb+v5Wfck+OPY5B+5GpPbOuJnB8yhgXATupu7gAQPOw
8Ra06efMogS1Sny+TPyQbyqWSz3gNfZfmqtfAUdBCWDbQuQeMZa4UYQG65MrlL1oEF38NWQhZV0G
8TzTRF0pqgw0Na4NVL11M5eXOA4APxHD3+IR2zjJAqw1L7MXHhXVRGVPbFmsjOvzW0MG3/PbubJO
ncMeVkGqd2KJ6ShmzBvCctx53ivKzt2ZIorh+3G2RHu2GjzMo1RdOwOC2PLtOaHFCP/wpTAFrz5L
vyDF7KXqPFgl9FC4lkc+4mXDh7dcqviAv/AH3c21NW/z5DWtyg40ePObDdeW2h2qRPPCzp9VF+P9
rfOItF37Ot7NicUOXi2k4BKFLiUEDPgNJCYjB1tb0AiIW1s3vcmKe/NGPlNU7IJRWZqcUpAF8t5D
44mGaZT1VLdV495FrImo995CWLiksfWR1c57jzBe5lu0Jn7TZrbPzwK6AKWNSHTnHKQJSHcWm0Wm
7YIrkSzryK8T//tZ1msb/j1TceLjMpxCpYysLDJU2DOE1x6CzEl005fHyxKe7ZhFORCY4f6Lv50R
YPV+K/ye2JwG4G8Vd8NhbwPfd/SkcORtk40qgK26ms+r9Ig7U3/cv/EyfJpU+Zc2iLvdpD7S1Pi/
N34N2IuWCmhBjbU3IN/5cspZdiUQLoyB6eJRk4+ZOj8khMQalSBxs5+u1cIZtJuQdwiayA7Gkxp2
cI0Vg6XTLEDXk233jdQ8JI7wovdv7i25aZhhvNAdR9Tmk8ENSCIIQMr1MfUclVL2npeC8mIf33DN
setGXNxp6+dk6whY92XMbR0WFEmjvtfHOcETqlxSnU5TSSb/CyNCmMcWQXmC/tLEw0wUaeWUhcOU
NpGdqoJdllyEavaU6cxqQRCNMfgGV8Y0WLKAipZnPZpps5c3pNtPpbd6WxMEt8eyJlK59yMtzCUa
ovukkLLVSFSoGKzHOuZIj6Piah7GV3wQ0nQi3h8hjay1c4PdR0EifPrPUKNd0lz06hgCQeIwSeSC
S33TrOSAIqD9Hgmq9igNmBN0nkRS1DP+2VpCNCcLPazYGpmVciItE5P6nmlYK+KQgDMepdyO/ipj
NuQ4TDEXKpK1QibceVde4tF2XWqhrPqXPoM3c5wfgwya57/rCl0PJ78x0nv4KQZ5r0nSBKhxKEEj
S/ylx5Pr4pSAaaBUNpt5lFNd8bACD/ATMX0dmUW2mhFXIiTbZll+28xC5Xuu/cqPPfhpgArNzODZ
NtFfCDSvmkMmP3X/YMQAYtJh0QzZOKxQSrUoWcYSPvIG+ATPBQUu7QrqyE/gLFSAVIKh2jkLKeU6
qMvJoJ2ImHoIAGAFX4jfYWgi1NvTxThaUKKYl2hSb9KEHDREdoSbhZb81r5O8XIWjueSeH2HdMmR
Ycw5a0Y3mshLirOaQ3qascb/p+qsFL5mTrUqWtrPKEaV3W1R5yXW1CtrHZ3QWlTgmQBL0vucEpxE
96NptC3ko7FpWpXQprTCWD094yY3mLe0fyWDur60Ua1d0dKcN0n+/ujcKieHe9jeZB4vNAiDWsfy
bdOIqBnZPEezhZcQrJXifQQZvOLfebeuQZ4+J3PUrjp53Rzu3ib/40PTk/xF5t8OQ5a2q+N/Rg+m
GlgPUWmowuEaLNJ7ij6W/gzGUIQPfdoXD7p+b2RMnfHWN1AsixXGledyV6U062aBlPm+LS7uI/Pm
rgr7aEX3x573hQ51o4o9D9KKMBZUY4mRFp2kVsjH2mVZg6Y4KBbHaSkq2+VgXegmxukminp5sKXb
4BoeUaGJ1RE0N6iJqh5YGbpuH3ec61S+1ungYSwIoYmyLwA6WZxncxoq4WygnSdVpAooEEg/zW3x
aV3WsYzRhDochVQ2YBFgi2UddZgHJ7q2LdOG0yEDysRHUKxjO9m2RSoitjJ8HonRhfsCH9NSDXjw
CfhO5nt9ySFmQI6D1k4NYfSnjnNvcE4Guo2RdwJlNOnmRXcmeuxqiIz+4cfmV9N76WdqAa9SRYQw
ZpubJ7+YCppCQpji4+gspgli1OS8Andlvi6cZzCumaRA3OcvsRU7WLPONuTWhBBCOptPtOJSDdpN
w8ccSH/OBdY5TTD+y2wp0ZTpRMUVjpixl0QVDjba3STsgnUVLsQ2+GEItg+7bzG3QLStI58Rgdsp
cJLi8IXF+s1UUiQ2miUtAmRlzl5VOTe/jTBDO4X8vcDlVSHNnZxi7ezgq01U7xYPucsImtGjlduU
UDNengFcAHNSLLqfhe8Gd2xBBwbFUIVCsFH/+PTGkxlATdCVgzET+TfgIqJsFQuzBXeUIDhI/B93
y/qOrXCHEArQY1npamxj218V10gskmWzjA5Q94ScN8ZIysGsVMNn7CEltW8XeFDZm9am8xFHyvwW
d+qEfKf+TwakBrHDa2QvjUIxDEg4bIMWuQlULhmvpb50ZF3tF2G6amuPzxe8aQEeU4BgpEDnOvmA
Vsc7OlHfiuztNr+IRTuZkC4yPKFse/waF4Fl03HOm5rBX8DbZ1fb8o9Ui8VpTAsvyp9hK9x9dxOr
Qmcv2rdIkhtpNV5NHK5iOAWPrCnzGEkXQOv3oCH/OwMlLNdanz4SmjabGHIcrafCrzbvXwazpotb
QvcVQA0H+/iFkz5aF9xZuuciIOnmipCO/vBjcqjJdgPpAZQcCjS8Kf4y7pJRy37fd0y9mkv56odM
HbHo7CTGqWEOdNKXsahQNF9EIjtTFLbPjWNj1NvTRlmX43fxinkKQoCClbAtxUPzIaaXR9B2L5DH
WjEKdisQD+m/fRuoYBl9YuybTu3k4e6B8O470iN5ACoeO7RKDp5wNPqeQ7+IMg/raOLacxMtC0+S
UID5EhfFU+Qso13AiBl3lPrrXttq0K7EdibaWSxV5FLPZnnypaImVFzopxEnlYpS60x/aDs/kHD3
EnMEI6yX/8TGaqymT3XMGJegtqBMXpz319Z0ebU9hn31YQaIg1Qt5qpyCvwfh8RYFH8cJU7P4cpY
dLJ2YtzeyPlxgA/gJkjZccEBv0jEEtuUtox0Z0AEtLd+wMPIsaf72FSdRp5CPKcQwTBI46OQaJsn
eNnV06B1kbS70EMUbiOySb8ohymQ/nc34aj/KCieyP+knZS1Hy/DQuLChODbBOILqDuSkxCbQ2sJ
v9ciF7PDNx7v0BeR9ugVTaRu2HoIFUGpdaRkdbYAaRNgQE0a4VpDAo1AuUpRbyz8YbTSwOKKOoku
istCiT0/ZR3aVH/5qwW3iIhHlEO1cewYUug4FlkP7VOWrQHrvPW+wQgJoJhxLaSdHgZve4LBSLrx
gZ80QN9iFVe1AJt69F0+Imn0pzXr74mJuow6RTZVerO5tTgpu7SkeJ/Rlja0mZkRcssPsJjCkjll
rWFNsnlbE1f3rUeu9KMyuiNIJmluS+cyjMI23QOZz0/RmyDFpLAhgllbak9cgGICJuXgKgiE6dQ/
UbL4JzcofuyMGkP5Efd5RhW8UcyVT14Wh5WhvkP/hXr0hfq1E0ucsfxCn6mK8f8l7vT1yiUJr+eG
nh+02xw9rhm7PE6hPilXNcaVu9Zs78ZEN+nN0AUWKGAwsQAYMmJLOM+efgCL6gNmAO5MiONYkRCf
Y2VVEaRt/IbCbTwrjv5JSjO13357VHX2lOxYfrjPOYAaLwONAdD90pWtesrQl86v6NSwoMAhsBaI
kA/79Uwd4/fEt8U9jzrTO3GnQ3iTlpSM6UOh+9G7OcYcvmh7wC0LoaCX6hvuJ+31EBnublyPmxv1
S59wIBrgF/Rif6MCUjxxtWrcEqiX33H6zBUnWajSZOnMu65N4YCukiNRTEvdlm7Vb8bZwP6mE8Ry
bCSWYSwcZAU9FUWuBFXQuJ8lL85KbmsnUufD5jfE4fN0AK6cF59cwqXAVF2oozbGwIJbUSt6rC9z
hZ8a+6FNcxy1Xn15WvsHTgM26GikOE6VSZH3kqrMhqHChloCPUw7C19ogkUWz+e+5buH8rFkyJz7
jPV6n7hcSdE0e6vBejI25R+KWz5Hz4Z/HzARItEcUDTqVxiTyKtPuWgJnr73kbIuUm6teDb+BIUY
OL7mxlD3Y+8bJH7QlYcQKTI+0pAN8Ym84BbmixxsOJsySe8hCULi8CnN7y8Lf1REwxBM6ao+6SoQ
0687ae+sL57xTK0tjJBG1JouvpSC+b1ievKAiyHH7rpzrgUG5CyeVK8ox69jTOknunZftaC3TZeP
4eUhekBp1IEo0iytvmgdxx1jiDGiv2C9bVnL8r9iNRwoq9fLRpRuxeJeijeiIF8aEHK3oc6WQnvN
Gt447/FoY2ejFSRXn7Od4/0vgKHxBZgTa+qlcCGtbtqGkz0tT9sXSSz/CrOS/zlOs7qvGNVMuBST
YCor2FlDWsIBqy3FCkHFfq1dCIKxhvTDDs3NLbT/c27MvLoXJOXU1JytAiKJX6k6hypqLmLleQVl
92UJb136JvwOYyGYhXkek5iXRnJHhxUMyMP2bWer60uKjU3uEnjcpT9hPsSFTlERb/4ivkQ1xZKt
cHGlA9UUveaUQqtZDx1H8xb7NTZajK2U2ohZI2nk5n6rWeCX4jCQKM+9rqOlRsUIrGq5W+lXUwwB
8ysIItt3JBSioWWoN8CucnB0x703AYd5OtjmL1IRExajjMANzlIhW3LiaxOCxwlpybaXsnFgw9aI
D4kLISvychShHTEYLzcF5vBMXFXtiyIUoF8s8OJGUSgvaJriXBXQ75Lmwgw3jPoqS1nhwknw2iPb
HFZP1tfxsK3IkzBQ/gbeh1vlPD9YVHJI8w/7s5BrXdjTvoTd1tibK723VnL1fha01iyKkJO4Eiqy
RtnkmNsfNx0EqIa85CEfGmI87vXyBpeZ/4hBJKX4mxHHwnOegc7xELWa+rg6PeDfatoupJBJ9wOC
RUWCTmMoxqHJam7pV9QVg2woQ+TzdVJdbSnAGltXSZ7udElL2FmRtTT3InaEw4z/bPzmbOqYmgek
6jJF/3Yvcm+7vpLoMOLNW2+yg0CFABfgR8Ljm0/UKtu4tSYwQgUOzS17KfVXvwtrrz9f0WbgX3Xo
/xa3N33vE1H6Sf6ZCQx32FG4bswhY6b3xbbJ5j6h/PrV2QMIraLSnlyMN2K9ZVP9mkMS3PWyhUYu
8ZLHVf8LOK7Feavi3/kBxVZbxdqWVqTMk0Ul5k9ObxcGnkEdiRWNDkVazPRv0gNfLBwG7iYGB4BY
RXWDJnJCoHs6uCKJTkT6dmikyCYlyRFUFQ66zGlnGIZWMwJqZVl1LK/7jSMjeiTSiazjr8R8lpEk
Z87c+MfxUHvQ5fv3CsXa/LO0BytJsayDDXzy90Kv7Ycb/f+Tmza2WXVNziqH/hzXR+IQuvH9aGNJ
BbUOt8sdcPajfdgSCvnyu/4qxmjKTQKo+DSYIercUDVkhu3LXAmWE4XeHHq+Qs4Kg8qSGJko6laV
/OS2tZ5sg1t57KznafwsQcu0zfcVrTinTmLAS9ThCaq97HSINUmVMG310OFo1MYTyaKQiKRMbNy6
2qgag9gew8lbO7eY3BZC6f8NPFF3KNP960g6DWWhRNs2uFM4uQ1N3md/WCTub6fj4yglD64N9SwG
Kn2GCOnbk+ACM5bo1CnKeFUNCGBIhpoRaIRlUqnyGJYDQWr2Whn2BSV2xW9k6QVtHAkXonT1j/gd
4EH/O8BI7BzGwzea+ghLx2SFGOZZLxGc/cXyTv4EO+X3FQbO18LndAqByPpX2n08B7oRvCPeTdaB
icXKMhK6lWo8bMCdGhLFDN9Kxn4Mml0KaTQa55mHkPJxzucJvzQZqPLdKgGt9RAxv54Nm9BCGoPG
xBlwUg66ysbfVLDkoOINDTJH6Su46AhcLSwGddF6WvOwkrNvdl5fpa5uM3ejp1z0yt6TPd3O1S+x
tXB63ELiFP1rwXj0GRaCnmvKCLZHK9RkttCQR4U1ISe4y2km6eRWwApNUZXXE5f/DHcFLwWs3Jl5
uKtXfOsM3RbsMXuBwvqSLohLcocYB/uRi/3prSHLZHPw4sJK/RFNSgwJ8YLRfbDcOGU1bon1AHu/
DdZq2AAqby9x8jFys3OwC2LuVYnecxVwet+uNch5YzhYgDNXZORPkQOpGPmRrdmKlz6ZBq5+k/h0
Z5F/2tyE9Q+bmLn9NRUT3TPhSyoSgwPURnFAnzogXr+ZeOMklYz8xluu7kWec0bjZh4ivyBhNbqB
jfms7xGXfWuRXsY4/mL6mEgUo4BXa4Me5f4TN88lQnZuzyFDtRH3j9hXvWIAgpBewq1nYrNq6b0V
iZ+Rq7PDrLf39IgzwbGilPkyHn3BN0UYIwgh9a8f/1QxN6hPRZ8n1V/cJy63ZQaIrpLyikrApzdm
auSug9Y6d6Zu1+cJHG+hcGTmMK38OTKzkdUKB/r5EebfQox/VUsafiNAnNSwLSM/461Zv4aOnMwY
O/WLGUN/X3ZBrvd3NL7wyueg7pu2f6QDMKHam0ZWrnZkwAAllD03r71lciXZeZm+iX08dYqDRZtd
somo3rJs+scBh1BvijQuPr9Cgo8J1/5sVe2HunAnrzZDblaEfmnPck4+QGeKkE+OUAr6ji7NLLuL
5/dc0BtsAwEbo7asvlb0K71Rsn74hc1Z3gCw2mcbYmKp5P8oNir3YRPuo2E9/hfhBcTno9LUHh5i
tmb+dNLhSfis1Xngj4uPcllnKkQmaqYtpcfp4RcyQUBWrO3ayyuBZ2nvXoDSTFyc0bt34npGv9ae
LcOALt34lVUhriMnAt9C+ZWVII/WDtE13Gtpv4BjV76/I1r0Y+YWbuPzLeiPalMi3z5fasgTcCvn
+WeFXz2ZffIqctTNjEHban+1HxVRBE3uPR2XCBdWtnhE0C5rlWRHNgQAEeY9BGO+O9lQ5+AUsKWz
7LTuIKInonCXHzemEm9b4arpgd7sVIu2j1Zh4/OSGg5LAsS76SRi/FXFfI8Xl8CYDqmFu5xWs43s
T0Bl3G5l0RU9/wbwcyhmmGma3vt0/h3/v70Bw7tu4gtUODDyjkrErDfjKCYXA4ecLxv+75VURLVD
T8uuyO4CODp9UF73jnU4wYDgRuruBeXAQCJ+vhCLYnt9rR6idSZzHSyNL2xybEbfU/4nOrT4Sadb
61dFSd86+wWJY5FhwCvoxdxko3CmYIU68praZj5zp372AY7uud0AVyeWEgC/4/Ol2kCZuzvECUho
a0mJe1t8WbCzOtFTHKjdaRfNgjGWS74vtiq3kQxAdZQfeH99wk9TVPtKs0gKPcZRjOpJV0vtCqds
bfgGTTlxjm/JxxQXo3wkrMeAdlJ0eNOIZEX2oPFd4+aiiCZSxSP3d6ljWc/xODv/zN7ElEMpKnUN
5upjrRzhfHKWD3JfWlK8PPUV4dbJnjalAJQJHkhk22bznc1Q4kPQyUBV+g3UuR2CAalFlVWsiibv
+6kq5TzQlxa2mXbb+CNt3V9/tLxYUjAY+JejHn1vBILnf18KkP6/WizPDtS3YG+NvEFd1eWwyJIQ
Okb4jQrIrVBrEC2idS2rPlW8A/ncBGkmzgcpevJRfrcMxhHropuLHaoosUBa2aKYzLRAIYtaaDGA
rgXdITeV6Npd5gpr2nu2L+knv3SfXL3wBmacLSEIIccUmLnIG61W57R0VoILsuYKH3EyvRV3YfN/
DHA24NiYr2sat2MfR4yPUxKm6DBsieTgknXt9AM694o8OKVDjuxmaLNmT6wpj6pPcA4u49aaHdTr
FswUr959Re4TyN5AVtj0ttTzddlfz9e+uFM1QgkxrjrRZTO5KGAIQP+uBkCgdvqn9cFgDONJjv33
K+FwYkRJGul3/xTnGxYtWUmPCcT1rY4UVveOY7QNle540cj3NMMT9e+Ap02bx/4X8dG7M4raZJfg
2nI4Gr7WgPGpdJez/7T0RcOgvcGJMfzhRaLqWVfu480zAynlXQEONbn4UTp6WT1OhIE1LEVLpQ/r
9BfEmRuY78Py1sEHi9uHZU2w0Cmkrc6/HP06o0ULre2UTDEcJQshNcRhXKEtTSsz3I8NqLrGkuP6
GkDIQTYNozAp/8mDD7kTAtRRTQNkL4uNwBFYspXlFhdFoFQQI2ill/LRtckooeouRlHu1HC1Jw9R
UhSgYbttIy7izW4YtHz+Z+uDQAphKjkjllf9jG4rRd7HQJglezW3H0Gq9lcGdtv0G/wUSuoQ//h5
4sooN/tUc1PtYrFZmkLoBJTAQgk/OoldYSvkRZPUvOwREB5VhOIt90v+YAhjp1ZwooB7Viu8bomv
al602gBH4UcgyFn74B1Rduc5XyoubmCPnjGi6SIcxP4ewDUvLjOMAUcSFRYhe6Dwd6+yxKiCtwfC
sZ51wptWKEYGatucGytwF1s1lOlxVPnCqx+QID/m0Qqh+wp5ZlnaSo7LbF7Wp4Bjy3Knj+GMd2Qt
t2ug6/enPavnQWASJIWeMjAB4VwIQp4uInsu+91HlOK/rh3qJh7B7r9kbc89EwzANSmhEmIpQ0qI
xa9h4DlysXd/DTXstr5zY9F/xQnO02xV+ScJXb5HEi6qK+Md60bLq6UOJURWsfoJ349NxI3437mK
r60FTYQNr6pgettQQKxUvEUdqW7U6xGLMVBLwpTtBkgd3gSsHq2t+aUrxWz5HjUY28yYpfNgBSr6
zPKBIvTV02zdZsygZ0iQnMO/RSoSJMGzF8h/fTTpHRrT18k3JI+zOzkOF7QgEYqyK5Wd6MQfzK/1
sy6Ot1X9vp8Qk4Ef9xwflaSHmd4IE3IGXjQHeWqNlgfwWUyC4h4v77SD6KGme/OxwkEMGu/uIojR
QxyYh1lVsufKXnOfla/0nuPC42K7HyYk9NGfhN7htXDZh9qlZNf5psyaMo/DYVEPCP1hd2xjeRJo
xEhMZAOwhsSvwoaN1C+mDP7j0BkhApL2ybnMHX+kbTuJM3351vZU0WSIigeUkdkuvMI04cvyhkx/
IX3fH7JOkL4pv+EpWlmoLs3NCh1fiTos4yHALn3JP/eo8LdkqOCPJq5UtW0VZYHY4Ob4QYNZjYsw
HMAzhPSH7CErABmq5NBKJKgU4LpTKcdQA0XR88R4sQd2n/MrVIil9tLd0iwrygmBVPefkkt6N6Hu
JAU3pwCWsDxChJswlUQiOoC+u3QOvHDQk0DPt6qqzBHk44J11L6LuE54MuN9oyb/SbDhep1JpFpu
4TtL0LN72dfRClYdJpdzgo+WzNOpdYRS8fhry9GKhKEJ57lo0qh8d9zaey9v5yNLzZ7H8IdfzHJl
RZaARN99tv2e57IpBxJ1BXFc4Z9zgX36KM6itYoeO2UwbyN2eDPE4SfVmn7DNPweNF3Sz7XAzxq+
hKM1FS5rWE33IS4LfivHqYM2228qHe+eE/R9D0VTTloCGh5FV3knslBFjLSXnKVAaEbLGzgLjuU4
XerRL6FJsl6RtxXMYeOnWDS0GH5Z1z+USGP5dzEPZGzBC67BW71DjeRPVsY8hJwnDQw4641ktlOp
wHD8EhTR68v3D8yGiKBHPdCKZQxWzN0n3W/AONNQwj/5kL/4CVH72PN4B2s080PILzRgpB4oC6Hu
Zmu9oTQHkBmO8TLYEzKppRScNxCN7OzX6DCdJhP8+BTjpyMtruVKg7DDBZsO1trYTl4jaH59tQ9k
8qrPcF8o9wajGgFWeeYJT1XN1W1hnOE2HbsyC/AMSpee+vxvMdruPZdkPTW8uXGHiyvA637yy94y
5zbcX1Rr75MGA7QKyfk3Pyj6bv1yLoPaRnWE42B9hMPymnVuZ3CazIjGyTFJTC+V4DYm1sdqeETG
VBCzEtFYp3Lj7hFWBrFojWY+w+p8YdKFmUQUO28Ofx1FNowI2RsSkH4Fx2zTjU3E3tMgcnyYoCDw
ydURgAb0CxRY3LrVYuuQitkxs5EsZTxoD5GNea/DZ2AitNeU1xJDt4P1BYDpJR7I6eWyZPQ18EtB
ymQMInwzCLxq6B0rDksE6/72MFR30lJSsNK5NohGHLbJfqQDHGyGfJT5px+t1rxNMQmBwz/O0Uv3
tAPlXlWhUy2nm8euEwyJtfMqPo6xhv4qsBqc5geOEAYvzC+Rmxjm5YJv6XmdL0EGsbAMR+x6Kymt
cyzYtYaByNqYCbshcXssC4mchtTU3YWYca3mt5oJv2hr96vypuDqqgScfJE8KSSZNutku5Vf4lg8
IkhYvwyYIOlMDrR5dW0NqASwQCrvpPw7y0BR+fRw/DEEmSgNNXsLN+7jNyS5G0Oh81rpE3eiMCyh
7aURQ4wlBrl6AmGAMpHt5XyAnnIizegOwXktCp1O9cA1V/IQuelZhoAc1+zb4BjuqUI/XD3U252/
Fq7RsrVUYg6lSRZ8sy5fk/nilbScHn9/TPnNMaYDidkvYCREvf1cCgV4GXhJTISwB9IbwLbB+Ry/
iw5+v9fTpEBJ96dwT3cTTJr7iZjbBQ5mMt0qpbe1nLR19INlvIYuCxHIh7gUXk7Fxd6/W8J/Jeg9
SR/DiSxg9qR7OgpcW6xmEB7dhZXfKFeyjkyJ9Bu5xDzfrIXo9im3LcsoF6qGyMn3mW6UAuMf49Ck
yBiCVSJHdBucx8nHLTHdIxh4DFUiLOGIq4BxznlkvZEtLK5m4SMa8+7QTIxPGJm4b4QNhjQj+KYa
9RdH2X8y4NoHfXg15lTJrUUPC8yUSwxa1l8SYlFXyttV17gg4WYv11v2o352lq/xjMcFP/uWaSgr
DxqlMyfJ+1fpnVNkHY/ybiAwsBIqjgSSdI5TbHYjc8PiS4AnXfFPH73E6ICy5vU03mvvKIlPcJvn
/9Y+aMizXVDyE52RLAYN291dIzqs/hmUBK4n+DXLISP4vcb4KyL2NBvtrk+lS/L2YUQpMAr4cCcP
y6U9CKdatZZ9YPUyiQX6siBWkaU0X+6hdX1jUqAFlq5epsE+VIKj5skow5A3o0NqY9WMfvYGPW+t
GKJbaBvL88g2D4VhxBwtKCYFE2W+kRRJ2tnJEUcys7+0d3ExEN3MlohHzGX5tAPsV8zo/vPYK4ll
hHi1gohYkhwa8PgDAau8W5KrGLOQfaA0d9XEHDbQKhoPqQLYfiScLP2XBsPPWkM4ev4eMQYkwzgr
J7UXvP4PhWNAfbgJvF8kCGS2uU5kNQ8EKyRoiX+oBNBoGg7Yoyze9PG4cfyQbezxuphkweuS9CW7
O/Qx9eLOn5Gb4O6wdIL+L8B/gIH/7e+4CnYvfl5WnLHr60VWuqWR1mYC/gQxnZRNtt706nrdRJf1
yUIpLGeIRlGkclG0INIswBpUvJZxQZO2b/5x3MKXdcbinVWicKAIWInAPuCEnfEnuHZ5acxmcrZz
IW7RRlzzC4qAaocfhCOwWP4PdIYp8YNPSIZdvbw8haSsh/goF/RJf9e69jq1X27/ELPlWmMlUgiO
N2lbMwwfLU0L88mMVdeZDN7XjzlrhzM8Tx4UU2ySCPUyqCOnWamZ4SD2kFBt9hWoPFb4Dm+bpUxI
DI0py0figaSSKeVliqrhFiMfGZWDR1XN3FX/v6ut1aZcNRVHcmWiOtXZe3l/j68haSlGevOiT6lv
jjtZ0jq2gS1lmI0fxF2Qk0EIXQ/N2wVnz6RJffneMbmYIjLUbG5Wxyls2gaVhrh78ZkxhmxBE708
w9xPjr7dcskMxjKyb4koz2VEB9FzkFh1oXqrT+l785Iy8deZr0dJUBhktkOVLegLQXHHw9G+etCg
O6F6Hpqa9KqlV5RGyDWRku4Cwq36P4ul122ntePuTKSYOvKFvXEfX/HoUC6GMxm4mfWepU8psR80
YeALXA4NciIxBaOW2m2lXh8QYy33CQn2DiAFXWuOz4vKsN6x8nI2oD7r07vLmnmSc60lp324CNf2
LnABEwo1K/UIVJwmfLu+eWZenYZf0YdOue6T4L/zujYnSlbZV0AWb1VFLVy56hmgS7m28Bc1KODt
xWscKaEnL+TBaohZXJdzH7uHXaD7+42uBAPylRRcv5EIRl3BAqlMBiz8l1eSx1zsY+/tjDXPhMhN
/2W38TIX/QAtZ8BdYN7MAL2EVsnh65L9Q1o2gcaFzd+1abcxWR4nRMOun4nCqPXocT/vZf705N6E
9LWWK7xHTGgN6Vj0f59YS+WrqMwCI+Zp3ccGJ3UE+XAlB8tMuOhTjHJMoq8bcxQXh4Y6Ob+sJmVG
8YsnxHXwJ5bdBwsYfHt2Sgye69BuE0gom/0cm6VECfiBraZiygamFLsGAxQ+8B43erysVPHF4F36
mlBblM53tFGloqdvxKCf/i86t6DOJG/AZemy55mjjUmfYIWeJo67ewVLwF5v/ybrTFW1FeL7e01f
ip1xwdUMXic+1aTa1VfUtm/uQTnI7+dOLnQY1Lvs22IaF7YXsOi3BnRnBUeLV8sHwO6E/e5Jso6/
uHjOzh39BTpzZ1SnoXbW84skQQmaSUbjeFuF/0rb+EEk/OvZoJ2VhAnWFY8eJ6zMIJeMZ5UGX/oS
RzyfZWDXiJ6wJN73QG8/RH49BJpD8gpj0LGJ+f0UZu39L7s2s1osARtwBFBfJ+x+KQ+8pllq6Hps
3qTcsVbj8lV+qJYTelwjtjGDbRpML3lWg4gQMunoKFoJ3pg/poEAGKQifw7Bmgs0wUdr2yc7/eRB
8KB/gRCrfE22o0nwORXw8hKMi4fIpdbRQAleughmT0teIyVHFWrgd/FQB1cJfS3CgiPIZbs5O//S
SuCFwJK0qU8Bt/aV1nx+GWgdfUWfeiKYR7+wrb5PqwJqV1Sblnfxxqj/VG9A64TKl/QL3c5ReweG
22dgkBdBTk9sGLPzmdgQw2iJXPsJHLsL+vd1J64EyCfiIUZugaAZEIXY7gAzKOJys+AdXIkCMpcD
afxTpa3xQywRPSSXJgkZ5jRr4Ym4MnFR2pZquTRQPS/ZPLguxG58Iu97UGbHwIGl1JnMhoKTx1FW
zNG4pov/OsDr7V5cgBOACX9kFw8aoM3+mTjeqmQeai9aiMZIkl+RmX3HaWyIBBYyxoHJ/RpcnX/2
lvrBYwJZiYCAZ/PSBK5YcPSJUfVP5LN6Sd23I+OmLsQgU18zxQw7X6sKA9jru6UKh8uDbg+UV34o
BuWwjolsiUxAVg8ZrHdRyCh4ivKRlfcum7A/tyW7+YRdgiYFiLbzdguwchpMaSKPplexTIfy8NZH
jc8Nq/Xc0Jn83f4saHmImLoUDqqqoBdc8BH4nH4kvs4ZxpY50guR5XdKewuFDu8fG/kS1wU/mZr8
izdpUPZdPR/RvVyJ6g3yahRiFoJ8slPxftp6HepceOnud9BQf5uJqfqxwN+RQgJC43nnl1ZBGvzr
Bvaa24R00aysbo2qmvwuW6YlzCEa4Qu05lWyBGkGDq9hQNwaYFalCqNy1rcMhch/6+kEkfVAiEc7
xBau/3cXJHtzUM6xgl7ImWB4xBnjiipV5nlpmsKMwRwbRwLN3418hjA/SLxVrxSWjlzSvaHiUaBr
RvyHFJ9Xeo4cDS4J969xDKHJpmekgcC1ld13rt0Dp2iLrzmaxDy/gTLjEcZcv3pUfNHjfe9r38wY
sZ3WbWTgIozlbALXkQ8tUTpXPnltUMP+p+dj+xesl900SL4FznNk2o9WX7dH/Nmb7FomIioq1Xr1
HHjI/r3kDejBNX6zfQ4A2BfFdG6Pcrx7xLVjnw/fItmnvz2O5/uPSRMOZQXTWDYm7pFCfT2hYZy0
1eDDevB6SHIlkb3S8drElZqic0g3nRa1OqwMXnHDSjaRxyfH0y7dIvCuOQKXsOy/bM/aMM8KQkLZ
sF7GeiHcgTAemoWy9nZ28vtbtgrzoDLzCUbyI/fRL/QrAgbEEztfQO0LXIhNP3pTqjWtTSMthd/f
XXQCtLctV8xxVzuy8wuMKuri/3krD4CCyfef50HnhnLz53jiuAgLhuzsnS/007mc+erjW/10L6/k
aiPGVQ5BEQLjsL+lHO0lad3xtLi8mTBc+hdwFsS/pHrN8hee8lwyNzncTjBm1pKMGvxxrCMHVOtx
eCxha81t5/qZS/XoxfP3uVypCOHdFckkZBZiPhkN+nuMnhGnE/+x78nLiMCP26dZ8XCSliljgesC
a9Ge2UaBOVXP7tB7X5dwzNjLzbft9KA4O56j+DiOZ9Kqu4BjwEpTQoUOcvtP2dYmGddrvGiW6Kh/
317NVPMoL0RSHyaH480GQE5HIRLjE5Wd3iolsAfNR3LAZNATavL4FsWBJ/GWFhzxZ1nzXthSuPh9
DuuKY5kF6iaIi9sqkM2WDKDGYwA2GpJbH5CubvFH7uMcO1Ovga3VWi7e610eAOW8/DEWIXXWHOQI
7/fEl8Q2aC/Zuo1vSxjb/bwaxBkY6YO/Em+JaqzKjQ0WNkoetozRyutqBCDBzX1IV2kD1ULk/Gfe
o7IS4ncaw7jm10VLc4WO9vNRbBEfKBUX9RIbpN8rYo+Vj/qA3ZglSa1hYtWVkLPIpnfi0byQJTRf
xJzXxxyE8Sd/apNxoPAjxxg0u1JsXblG050Rzv0UorrkA64EcCC+qr/TvKCe7in1nA44up1Aa0Eq
5vhX92wYJd0LOgoWUFj4d+0G67Hsf05oJyDgy5bsO0O9g9zCCuq/n3YJNlHrqvxRUnlPSr3f4zsj
mDv0LwwPzgrJeSdPpCVvVw0CCTCf811SWY2C77be1a1Gkbq0/bvqTIzVJwy+1bgl6euc/K6qak2M
KpL2GZVC4y7Jgn9/uydDIq/wZShmyHJ06mRGE89CzRRxy+nVw0JyGt6bcA/NmPvjmadKjbj+XHQ6
ZiuZvd9RYQFS4QuV3tReVUCHfn+Oz42Ca+ZAAaUgsyJDf7xSuQkj1+rSweF7nA89dGQFKyMiIQ0T
1mkNjLign04e7KvByd1dpR95rBvTGEmX9khZ2hgUDIuKa+9PRRIiob7hVqHcWlebWwmDarDBLyQK
HhHbIXyIv6+mC//2bCL0PIwoswka3ygYDuokPNcgRO94D/ZvjCmnC4nwoAYVDPkvsu0kEpodWnHf
2hxYR3uFTFuKstI0nitWXchnQvmnQQGgtFAUc8k3rNnf84RI9PMNod9Pg33lVwWU8HrNI5/v3dEg
uTPbPXvoFiGbtbQgdpp/B7i/oJ98/ASbZ2ENWFSK/GJbVgWXWlKgCG5HzAPNga9LL/RLl+ahxyyU
VsY11YXfliaWagDKNLtvmYoMN0D+uD1xl6g7JY2IDchgmwHNp5cEKj7m4/urHjEzlTWeU2j78FKm
jhn5I+WUlOoaF3/Ia69QFEygT4WMYA5RgYj+pNPdxrA8h2g+4bkoguIxo+fX0a8Ke7nfLTtpumGf
ZDyvUaAARdeMUFy3Gwnao/6O11yGEDbz0mOqn9fWQ7MqAkGIEz8vcekCc1Xxe5ERkJv/bzWZ0lnC
SK8YFdiT7sNV8cavMv31j9JByRK2SQCZX3Ic7Om51n+Nkfb0ZoyFUaLWekqpEBYkVV/AW3t5g+y1
T+oeY1uCV8fXmBIChhYkeNKh1Ak9qk5JUafLx0Pws9wBNiQtev4tkU4zBD4ggw6WSN6P411mU8j2
mkRh1o3u/hGmTtUGkLIP1s4GfTR4mXEct1/NcRfa71vChWv54geyYJ9TGv0GNb36CnNYDhlSN65c
JNB/9lDJb7SulVrwjfO+jWtc325p5WKEvWodlGIzv/qDUNso6+xibaIxAEX2E55i9QkcZjtvaI02
AHIQ7lbWVsFmNaJKpXUAvtr5/Zapi+rt78orWldRalg0jrgsImz3Zc49f+ezxGUPDlXUXZToeZSc
9KSjGE6cfxRrVMM/f5gl1inVz4nPwAL5qfEkcedXDVmHHuDJVcl8x6WGzFN5Z8WfvSPZ4jzGu+aV
zNdckSbYRGW3VRwnc/fpfHOJoEJl90ujzkUq1aZ9MdoPKmWkzVYDqu7LU5s5Txnq6uzFz+M74l7I
JbG6vy5BBaCgIWZjz/3Y1a5uruanhKYlWA5YjzDgNzUhuYK0sH6Dbkbo1Aoz4fB2kxYtOUiLkm/S
wodWjujXc1GDBVVS/cKs+iQf/ou+JIg+SQ6zlkDzn/Dmx4TSxaVnG6cE1Pq2SecSPgxH0Vc1gZ4h
IOVmIQkd5ZUTE+iEfZhZXqLxW9EH1xNQL+f+w8LM89Y8Y+NgsgT0gIYHY06SrrQG00y9s/rBMExE
sjcpWqrLjiJ9E/jd5l+hQu/iO2SZlKk1jWrm998u4uqlPyLiOudMPV0150gPIOVPWNJ6k3VxU2E8
tUY+AycHNc+NK0kx3Cm6W+at4oC3WZMW/nX1FNdL/tq8OtGRTFu2CUWM8ZGKo+Qr13aF0TRkM9jc
HWosNM7/BIjvHzQBg3XD/UZyCoEG07TQqUwI5k95Kai6aB1Q8tJWZsd93vzcj73De0TsxbLbMxrF
uHsa6wnqC+aceM70YMQ9yKQ+o5VXytst51V26ByzFmJ3u0Z+z8m9TLc740nwoaiQv20RfmTgE9dM
dPZE7PNlVb+UgkHFsCaIyPr7SwdjFSzsW2vha5uDOL1GEtNYVRfjLst0KKF94200kB0g2HJiXBvU
y1lz6Byz1lJYeM6I7VIPKAhrAz0AFLEiIMp8/MCAhzQM0P1PbhOyv3nNEj0wQMOalELO4zCvymnd
pxXw9MhGK5NvwH8fwY2WDxwGv0o4bALw6O2Gc3WMf38P7JNoONs5DCfeE/gdToo/gesbAHnOq56k
ozrsxt2SdAxPYmCPMd2xiedajJJsB2LLnrT1TNZPYp/arwvS/h4CPa4aPRDo6mQ1VSsg2OGiHnVb
9A2CetUESixJaEiGCPXgrjiWxQL7SirX0OiaeaMTPZywc/RF5RirYlXMe0usEGsGOKEZdFfVapKE
SxHYyj3IF0ITWHdc4x8M/L4w90sydMAeDaLXo4uRwiDqhbkGEr6YsPBoHvPopB3gnmEmLZTTP65O
zJMQUIkUA/NiF2G7khaCvjU0V/EQu6QkQLsBLxQ37E4LDXGBTg5GEXC1ugOqaSQEtS2kSy+Rv32M
0hxuA3GtVKtsJjXt9WJ5f0MqEshLjITyP42OXweizWtciMuCI+uDODjn2AY8RH6rJWtilgVmwbbG
T0oF4qZXT02Lo/Ecu438V1M8N/Z1ipnKBasg4USadVNEIxKDLvgNFaCwGTVwfeyXwkxP4noisKqT
Lbnpr0R1jZUeFquDI7vRJHZc9nBU8gMAMNE2MWWJZ36zJmALvT5VpbY02oHNKW2E08IBwsM4+v8s
m0VxdrRW+O6XXmjv82gfiJC5xwDw3ecRsrTeE6tsOtMJXosWQsn263z6xLLlOsAhe+Ie4Izb1wxE
iN+kJ3rM2VwuKIAogr1q3jrzyAgguGvafNcRVaepxgXGQcCYZRBzIxU8nBJNIS+MuHsltFRzqUp9
EBCjRHJVsnj3GNtQzZ8BQUTqbHPmn7KNXs0AG5K7WOeLZGNFQg1WpkBygfRUJNbFaxbXkeiUiqUR
axXFF8QhZUhv5UQZ4921oL2L5vcS5Aa4cFU5xWTYwYnYifGVtoU80K7YErbT6ccVXV/1LfBJkWL5
XX11q14Lklfk6F4hg62AnkTiPVD4jSKRZOKojT2ft+Fs+fNmoRRuaYeq84CWYaxXu825jOUaT5R+
pnWsL14GzP9b4mWWbkiw/9mUGfLHXnvFnA8qkiUj2FS9DfobIpOfAFLOMzhRuDP/IC8Vb4toS2Fz
0v/irl1JtfH2odvadGjLMW6vl1anHpCMGqVMWPSI4xbSJ/spYEJHv1P4gFYjY8/NKLFGkydIa2MC
lWbv7kgBtcrSHTRGdFRplzI1pVlnXNxZ51ugHeIVMFte1UTD+oIj94MpOsbd9M86wI1Poa2zj1z2
GdTqSDd7CP+td6gbW7iUO8e4Vaf+fKc2JTkqus3SGgx5yP0fU0q8+BznHkmT0U9kFQiIOtS5LRD8
/ncJdEs6oxBE+XhVm3v4KgufEL8Rm9csYHE2wUbfPqaoYGtjmuq3/XZVOZElwIb2SCpxkbmepej9
8XB8/clQG13fq8eqmVF7xwjgxzo8xWfuSxKUxobM3hIt1yn9P+WxP4aaziSXCi75KQJ/e/4q7NVt
Au3oI7HVeB41kpM5wbZiTjKyC6G4B+Wt55VVVTQLrQ+H4GrCUpIYSqpj62s704Q63iBgM1xUaEzQ
s0siAMBSKK/2WtY0jhDTuiSb5zTuLP1hE2wPLi1zAkTKtb+OG5PTA/ZSTlpm257UbRJKuXkePZ/Y
dB1w3xn1sz+4UKMCyqS9Up/fbEr1Bsq3jvbW8+Nji89DwQUsQV1FI/Bw8GqaqL18qqNNMUx9rfy/
OC9TJgIPs1NG2VEoqyW7YFAGk74CMJ4lv+ofJW6mxgg40zOJ5ZnL80uYraAXq68BMXDGpQrLajbM
hxG9O3AzSod0k1eyxjVYyjlZq37VVwCPW/duGk62cJm7MPLtrLaXDEAmtbvUxI5q5GMCYQVuXuFU
uR+yWpsJVPJO25z0mwsGKr5DTvKVMSNmHWT0HIEPcDO/vRSc44RH/WFVM6yMRgfMYDeuTLcVFEmj
n6e5GMFnZae4RiRYucYt4jg6YFnVWBK+yCZ/Cbje4b1Sf45n8hpGfOt7U3MkW+1mqGRhDsj90NY+
fAXnbw5TT8LKjFrY0/OxZzvWsR3JXJ1Z7ziy4ToxoB3riMDNan6t1wgprFxsiO9vzJkyq7XGO8UL
KghAnj8qxabz8aDduI0vimxo/lWQ/9b9dZQgrzue1sfwgue0QOdQZJ6mMgPbIUWojhiXk+weVoQC
i0oIRRnJhorlS7yLRvKma8IMjEaJnrjtVLW1NxALoDMXM+7zycq98+ADvCBAvYmj3YA1P62GhGHQ
ikvjC2FhlQjoxNZnhV6wj2dhsb0KYyQC9jPO9UxsNMLFQiLrIXfCgsIOVrPFPmXOnJpM/VaDzUQm
ItkjGseaq4LGkF1H4YdKWTmxoqlEmIApoN4z5+CuyFDeI5lEpgXr5ndjLgwZw24IGooz6HIY9vvy
6xPdOO7xpo225ddKsH1OU1s7QWVyVa0PGOw1gu2QHJFKo0nREp8D2C4Fs7KaZwOAFdy/ZUSP+5c1
fkK8dpgiaQk/Xuy1pI/kEQ0GYWu+u3yYgQm7j1hrRPw2c5IrNw0R+UON8gvEmUZu3Ai7ep+hYC8q
wtIAe9A8bCOdJUS8WbRERIaQ9x7XH9GBpjSuFkfF5lGEWmMex9r1StMIu5oGwmtiX/f3yllc18U2
eYNiVCvZufqMPmrlFRD/bGrfeKBx95igHx8ET0aDm4zYHExXOM/JT17nvqr1m3vUWW9ood/ai2zD
28Q6z6sopkzsslODr5Oc4VUsBD7voirtIb51QlPucad98+32oQTTOxP4x1oplJfNnU86Yr7As6WR
HC/OaE53g7i0CTtDXmiD/n8HkEmjtCDXDsLWo4b96S9yzqDERgGSmQoTuOycw3uafokH7OxQt2fW
+VPKyLxxa44QmpZCi7f1lnGqWV9ikQHgyRmspgvoiwalQmfOIZxOUe87EfG5v+o8fJ/Pdp95c+3g
KAVT0YGf8I06aT5YTcpagTfPp4rLNX5QqE9scj6qRpZYBjeDRJBKVUs7+0E7gjTH9PJJd7+EPQhL
UZt2+Y0FjfajyyYLmaEztKOBgdYvFB2pW94+Whw5ADIz36MnTwIp4QDvwc4W65ja4ptdAWosPz+r
kZiZZyJiPkmNfD3K3kpB5wUaEifGiGAG79ptPAx67RZduKLJl615Sdxl/jNx9mqqfgcyD9TkXPHg
7Fltxg5/kfpqj2m63WCR5NzaWUMb++XmvshpsG4MfG63LhHEceNCBYf+Zn7/7AjcanotrWs8Lzhi
BAZVI1bNbw/kh38Be16ghPJ0bqzZa9WaEqskzc8cFZtO007Q7ET6e7Ony/4zl1dK1fObpyPhmG5p
LdPr7kiy0AKBkhOo25glC1YINsXPpr54ofx3AXT7DWYRwav0cVkQqOH1SDyjQXyuZEULW5d7gb+N
s8q70YzxAdK4pqlQNsaY5ABC2tUAm0e9tQgtjWJP8rmlLSeat5QRUnuI5X8kK01pVl1tphQ5QVjw
hmFMz5bTpg+JeLoPUmJhTYBWmxMmVRL1Oo4wEIsrRD7Ko6NgcJaSFYgPTvsna7HdsuXlct/oy0O0
HHYarNRZ9yr4W8UgJIm3c2J1zYZcndEdhv9xsFisYJi1kXdnPb/Q311O2EylIkTAVRWAG3fY6m/M
StVqG3hqEKoj3O5e8MCpgCoFHhKmdhJU7zUGIzm6t0DSXi7oLwqTa+HrfsF2LWVM6NAaQZB5o+9W
Eq8Rly7IyRjIHl1KPcrjW+DzFQz6j9CmZWC0UplXJu3/oGQx9l61adestXy5QuEs3LrLvlJw1EYO
GuECj3nh3awmWAa1KCKPJMURA/bL5HDFngFZcRlifOp09iYXdl/EWGGoeJiXCPYXyIjdCFdcfJ0B
ib806wfw5fjtj6FGSJJwJamH0/caLOjuC80ZL2ZBXP16F2HTd60kM6dzSwMJYguBP5RPhuFFeMKl
KoxsKzXOr+qDlUUYM2W0H4bulCsb2rhX3LYHsYX6jEswYVKLDpltK3sXxdpmyTAWY90+ByzjL2Fg
4b0I69u1eMcwY24Zn8KzfOKM/INpCo5D2FkaKcJ+rBwJ6RbCNlrfcEciJkG1urdC6Xuh68fa5SUS
NCnOvxeLSBIRZIZkZ/hZ8tFQfjjdlMuKPuHyx5W5ZUE0sAmDnFbGXhPVSZaV7uBsWgF9N367dbsj
NQRHv4p8HFDOUE/WXBt7VM1XTUx0nJ6Xiex4Vj7l6Ch+rvg8v9dtpmdyzagoVz+Y86tMq9cOtG9a
Rn9+UN0Wa9VT7eT0imKHlcMFCHUt8JK8raTBWLfBZ3tcA5VQiM+FEYMzpedAj5mQ3fMYphmOo4e8
wI3dux74y733tKzf5quaZhnnPOoTKIcH+/WAn7Ek0qPuzmLMVM5ghEBSoM3lsKJrcIhPwaoIefpn
b+R4PDgLNkkBlO/PZGgcPj5pdH91PkClCJYBteCh1QaZrv1pyBgt3o5ePMlzftRdWbtk+rcSZ2CY
TK2re9VIBJtpUFshjkaSLSdRg8TEYwYZFaIm103X1v8gFYHGFj7FF4awrT5n97GwpPNByATlVF2S
auwxr31UV4QmbshmyxkFBDkyNS7uMYsU7UBaVrHHLx3/Lsp/nYPvR01pCz3CTOwflYIqV2y6EnjR
yobNdOyBqCtIqW03QkA8QjyabxmX9cM+CHU1KC/m3Gs9M2k407gI3KC/vzFnKc7qg0resL1LbSAy
DtfEH3IhqgoWJjSZ/7G9ivttHqLsPmkKHZKo8VCVDopi0XzKk3fbC40q+OQPMBS+Wmm1trmEDaEp
HJSKnTmw1LooTBv8huhMRfNYBPn/P2xKryQHMVDSU/8pK7TNJAQxI4jlSSMFk7KhRMCx3lj8G306
vsN0wt0JTW3QbJ8j35l27EjN7SDEGZl5cP6tgmzeJqc0yfgY91INHQ7BqlGmoX8t+Rw0nBaaqntt
i7KHd3JItZNYUrPxVGAs4iSAls8VDwcvMZGyN6+pEEG3gDU5qQv5lhjefYWxe2wgvZcv3VuVuaek
ip2qjw9FdNXyZ6BplhWHigQVYgy4Oiet4Z5h5B10NSqEZ/x2Doj+uzpVt3Sk6VLP+RapCfJKrT/B
JvELMBf9IYUjWXNi1i3WzdOGT2q1kQEDA7URaSITgQr6is3DvLBiUF/d/ApfRTvng8PjAXwKBkdU
b8Hv0q30BdVoAyOr6SD1MjGCSlS1eOXljBsq66jQt1hjtZIjO/SAOyUyRNbJyvElz11QVqNzT7rO
MV9cPKSkKvlHTGUApZHUoA7dSskr5fJQvOscjvRaurojNBvWHUaRsmCFKDzbKrfyKzDlv83v6Pf5
PknrFy2hl0ndqv8VRSI30QvDJl1q+csIQyVVqCkAI0bU53Ri5mk1IFS6lsO1kYl9Zn8abAAh5IdN
Ms3yYTyKMWqa2S8LSoYxaOlPsoc9Sav0K02iJd0/7zDcS54Cn15cfy6szVfEoTweA2Bu7nj2pzhx
V/zhXgNaOC6DQ6SB2u/qH0loZHXaG73FaGG8c5Z9WhGpoJYtfMjvxqydC8oEN8IYQryDiHVVaDKt
pyprroBpSWZuXFd7Ww2/50ctfyANcqWJS4TuK/CTyBk98nLXTG5zUw0EKdnLkUF4/+UKK5Ey+x4e
ezDbi/vNOfgBtWZOWuB+uR+SFfyHu9KHzCMpmEItjeE0WWPFKECXaLvR7E2weHqtosNKbzBih933
AXAv13FMYajwOT/+HfCdgXWn9dn2ffjAUiT1yHtn8899hNvEO+utudk/SxDxbI4UhtfdLluAa/kg
3NA7QfLmJmLODHGAHAEbgmDReO8UDOqFjd/et9FmWhv29TxNIJrrGvZxvnG2san4+0JOjggj35lW
3mb0bgFVp3tyXvtg4qmTBLlypL2eSdHMq8MoJR0Sc2AofSv7cF82d1802/t0mpWPK4fdZy/mh9lf
c9enhl4m85DTRQQ++SCeXMowy+gVR9fD+ol41JFthKzrlqL3EzbHBd7Jv2owzASBlcGnQ0fOkDR5
jLWWCl6gIaLcqucjV532WuX+n9LSNFsjNKGk0xkIM1y1m3l4xjdkeATn7TK/L5RZRCUHttKpltTA
EWI2GLX+iuJYN1QM1v8Aun+aDVgsTKZ3EkrFsgb97vFUr/WytqteEiI8tvUUoGeGbMDjRWEtqRcG
seyJzXIMQLFzMO6nW3Q8lE3L7WGIZvHmuv6cMKeubmwPi6Ydxj4RRsY5XorR0wjzMRR+mQmb4prc
wyW4gDo7FnUQhhUGZw1m7gvo1ASkha1Msw3wC4LAZ8gEnVEku90em89AXZ/aG+vtywzq7BLOa3bl
aCUUIghNO2RIljM2V1TX1m4cGdfkOecHtHtC9kRCY5XtJydhkpH1JXMW6F24tz8dgNlx3l76L6oF
fc/dQQjD6V1yTBgB28dKQp3yMh9DiSL5DlKm7cFXah68iQo+6U+gJzDAw07O6dt/SoeuKnxfCsQD
CgpobNGQ9j98gF4wUkZJyCed669FGMmjNz6Hvnq4Xj0Xj3Sh+nd2yleaj9vnPsMF13rBAJDqrM+e
/6XCvOpqCwWuXjxkby+vAx51oiyZY6uBVBF3ejFbMeeMXnDS09dsjX1f4E4P8wsedHWhzr3NPxJN
cUygY/nR7igx95Berf21OcA/uWLoYZ91IIWSDlFe5t4ngJjA3jLOP3Ho2upsIxPK48xMDcRLtqgE
o5jKMN1LjK11d1CwDzoRtlIgI8u6qwC9DUUs2xA3zvtgDyE8hUA6BeU0rIbzhmYHVzD2s7j43jfb
vRZFd6iTJ6/n/lrrCmiYWEK25/GtuEl1LtjIEXSG7UUK3MyUPGSVzcBhBmJYS+EbUYNPR2baOnzC
oK4+9OgyVJq3ZUrt3El5hr3IlRErDEG2biXPhzr92OT1TlQuPn/PgVWWBZ2Ov6gQ/VZxUljB5YMm
PQJiqx7t57mlGs8XI8hLpnucYSRZnGjZvHpNYzLW0futLX9jMsZAkgTwef3NZU8cN+iqIRMSk53K
0s41w3LqxbILOOzBlX3722VcG7CofVq6x3YALAXWZSd5wyvZdyHVsLpz/4fARGvBwgEi+oGBT3mR
F1szgApkYO6UqVOD9vUH3yzj/MUxbkauo4NDUhgI5jYwN4nAq1HZb/3lIpROHYtdjJZFbLs9GDWg
egVIr+VA6uqRUQiw8EaQYCZ3AX5puubHzoGUqbZnyzCb4t9rlCzKeWqLYwqXjwuIvaeH8SyL2kdC
pITSppfN6xOwoKHILUmLOySiKaYWNmTwMKCMcRVecNXnP7Ktuh9oe/oXuH6lPDle3gEyGehoV6ui
lhBera9LyMM/+P4CC8M+RxjCzlPw6HNwWmd/nmS/3LPg6z/il5TRCQu4fPc2d5v6CN/OdRbkLjNs
z3COEsy9CL1vySPNs5bHibfejuWPQVKZCqCoh4d2O3z9cogG9PsI7QzjWVwJnhjHR2gLtdHmoCQk
yIWX8BlMGjIvjFG7G2Hksc1p5nbiI601P+lZH/zKBS49NSyR5vyUQNRpF1fR9FAhauUrITW03BZa
MR9yA8YMu7Cb/NYNfoRPj/umhpfLNj1F8Xf2XIPtLxg52/nPjcPY+THp8OTB5Tz+Z5eIL8k2CL1c
PZdItvPwp5G1LMj5cbQ4bRQISVv5qOzHph67pL387WBG41NY1tOVZi7AwWkaTCbdOVygPGTX6ksF
g8YftFBC5T95/93fbIzfEAJ3PvSo1sVMq4KT6Ih42wl9crCKycjpw2mO6mgGjq+m09gioihrAV3a
bCMqawhfxHUypaJS+ALI25pY55T9z5JtyyiKQ10GFy5hj5LPd5WUBIiANIirNTpSrHZkWwe9a/tP
ogPBAzRGieALRdSGY4sFbljC3gn6cmhlIh5Ak7fBovHwDQEOdNR7XtzlV3iUg9X78scbWCHuZ2yY
sgHm6/0+SxG15UNc9GBRiJsCL5hX2IJl0ToJGb4i3aqBm2MKhdwq+M6nSzBDER3YKI5KHf8GcBXD
kXsOUoS/5JlkPmbJyM3gBaKtJ54zwiMz+/Z0CE3yth8rxyHhNjCZpNHT4+hAWVf9RrY0VRiVFo94
J4raaGf+eKhZVPDSP+WkUrtwCeF/81d80AzHArdRoOJC5y7MSKLSlUG3sbUAVt6SxbLfzIakA37H
1O0rOlRcR4s2BThuphvwGC4XP0B8CfRbuh0pewk9AvDeEg1tC1V2qU98mh48Xvi9SleAFyzLhSxe
4SPkmR7neF9DYPEfQVlQ1uoQ73b8Z5YGjUD4mJq6jMUapDHMU50x9vzy+WEmMoCSMK8oDFOlfLto
cpF9sXZbrsaWtOEVk82mCHqJqnwEa48Z2CQugexh2qaZiz/v+UBg+4n/UyVOy2yzeHdjyX1l7D4x
lPx5y4lnmnUg5Hf4i1AG2vVY8/iDBP1493zYXkZ6tH74DudG2DCiFR7DVzs+V1pkhDGC0nYfZghy
k4too9/3aMou3Toaa7SF3X489laitkVnjST3X0SCSwmjV5+dmFsxv6x2CRLleUConNQS6aPnZR3w
03ILbDsNPG+X+u6pWyWPtP1KPQivFtYPoI3MOi8/D6SHw8r03dRApkL1/+dQIT28wrSraxqMJzAo
AnJ3fl4VMtOA2dl2/Bn8c67XFN6IJDl6LubfsTItqNcuUBYmH3dHm760dIJNrVXbBkiTiCXCKi+q
vQUbD1IsDveRkj7pVLgGQATtMsBWAmXaJwYjq0TDbKVIdI3QVsM122tACz+/gpY2UCoC8CHuF4mi
Y1HevbBiT6nqITKMN2JiKX57iyFvzjF43Rzp8gZXrB5HIot4NVr2Z5hJZmtVGasO136S4dVgfvxh
GS+9X4NmTY5MwsHAX+IhlktDE/UzUQCqYkek2s/7cbeilBn764ai+nKKwZ0LpTgrukcJkFB8DbTs
HIY1qopSKjY/P4vd0L/Hj0EcKV2NEX0NgBb7ub2HafZkZbEmZHAnqY2qwxoRPvTnIS+MFIdjfzfT
nOa8sg+Epx9eB+UcsJFfi6MirjbVd7tcDwYf/E4mtNXrfgkGS4nVcdJvAsdEnkV+Q5YUGVuoXRct
7MzxJ/ZMASe0ad7wQSIQmPVscOJmEZI5ZjkSFT3m+vnVDM6TUNF11BIDG8uqLbah4IsaMUyIRZnC
EdASc4UJxMSKWBJjrg1QhKjo3m6ks9ZnTcE6CUtjyj0Cn++8FunGw1bBQ6nq3FhbHxKM4ttjpTLZ
3f0zmDszeWH+zMgSXw5/vCp9XGs0NmSrvPEJSnyieNzZPnbMWVMVUZpjLOChZ+BiIPfTwD7bDFIr
R2jFAdDkDXhTV85xNTGNg42Oyg7cJj1xYherUZopKgbjgAyF2nzMNFgvuF3me/zX68x8nDgGJ07q
ACjEq42Ja2aGzEiToR/jUbHNwT06FBt5D6765v6MXAaKRyzOH/vNxLZVRerP4hmZ4qwo16H0q344
faF++Qj4CZ+1Bd6os90i8lUanoErxFsPeRDn+5mbuzRCQIwgtP+lERtZSwr8/A1FDC/2PDmkwfdh
sQoTGB8ZveP1sSkXn7HJJwLTF+R9sdncl5a1eoOVJzF/ku99owGq3Nm5tP5M1IJmaI2HlCz/PwKP
cgOSINuIbcqtjdfkOTNudSnkeJNBv1klZV1xoy3d8wG0vIkSNgjCz/PgwqBACbNmsLCGPi8Mp6ck
qyNbr4Dk1sd8sBF86KOE7dE/F/MLApRG9EeQKQAn6Jx7y0F3sngkRLVag1W6JdXeRizpgj0HgQmJ
S17DCOyYNlNpXbK0hmnTkTZqJv0irjBnwnb0myEFie9CzbWpVjHfczL1nhHggCB/AFygIGwQgMfE
wWhng6Q2aeUZ475PFjfSQQ7+cK1rHkC/vlC+JPpt/SbrYQ3gUYqvddWEEoNuNzPat/TAdRdj+f+X
ZXl2sBeKw1ZWmzlGRDE/VEef0Njg58L2I3fmYI/tBU18o+cpxvr1x8dRwPzYMrec0kpjbzXI9ko/
mc03N//HNmkemqlH7KfkA0SoNCyvCXqXCR3w+7gBlcQsuoNd9S8X8UbMtGpn1Qm6hQjx/KPpaUhk
jMrKz3VP9iXw5cBQNGyuSovaB9c+4TDMLYkRVr+J8EPf02wGpJRStmR+AxYRUf6KeQtgBoZdkj22
jJG5qdHLft+lL2xagJrSUyfIh/3UES8Dys6LccVEcLHrsrzlxk6G5chZyA9tPGdNyUHKxcKFwc+m
lvhjNzBFggTsQ1qdvoXE7KpL3LPpSpxt5pRqpoXEDOP51p0dtsx/mdnwTWt/3lC85tsWqrenUV1X
V1y+o49RlJvAFDFdBvA0HhgPtjC9PLetE9FtBM2U7HHpAXoqmC5jTC1LeXlVXCShyMzR7asBcJ2Z
ynZIZMVtqvrMUpimcy7swK1rWxNCKcbGQnD5O3g5I9dEvQrCUaVB4rAgtKXpVInLM1mc9PsBfFYf
jWF43CoI94JNNizG+LvFdUyRE9rWV5TM3b1p+ATA33dK2ztzAWe1fnbGisTedkNrgOexWgfD86sp
Eb8UEKO+5n0/PIy7As9VJD/bsTlzOyYF8qUwAwOX6WO5z+LWbWGYIMcpjykLKsiURFODTJSQWSfj
f7K44tlaDgwaN2np/xtcXBtWhcGNvdI6shBemgu3TZCg4kJSMwLiFtgHx7aui6wnLE5zC5Eo7JWl
Rfox1rzQAqGT4bXU9zPk9mjcSLm7l1DFq7IwWFt3odwaWXZrjEeIolj2Vp8pMWJ6B3BKmUMPStm5
l6RkMStivmotBWT2TsZWag8M1c30s/WwtBg1yey1Nb5AB3n/FKUX5js+WIA1q2A7Hk+tlaBsKpJX
XTVpCoCIldgzF7gXROmKzleEzcwAARi0XBqU3c706XwTm2TfO4ApD2PA8VDWKVJqqQRqJelJeQW1
idT0A/UxYJgcGsnacpEvK3yKfmBbTIA7V16gP0InffNCPEPqkdxQ2QeoENGEn7CMRjlqyayKJ3up
qzqkkSBYkD6MxEkTdt2OGvtpMcRGABmbMAwpts6Fmw23EDyYSZACJSOvSsRP6LlGAdxf2Wmfj38L
X6Z3FM217TBHpF/CAtMPFZtx2gn+nrhKIsSRzHlMSpZb6wJZ9mhC/4BbCMGfFhQEtFFF6hNBAEjJ
QoUSFcTAs6ySbBF2FuHVdOmHYvvcIZTAkbdyOe2clU7+VpekiA9k9csoObXoFemQQFATRzi0CF4u
t397i24OGBHU8uxaNk41Uzqpb4/VTCk3N2g1MN2msIUEgKgBgWoTceEmR/YKJCYtttrLIuHWNXi2
qNk9q1NCh8HCbHhhQCUhudfMT+m4niqOTPCuNKEwu1PVwYOB2KkO7YZXGtR9YQq/h2b3fHc9Ft4l
FQA5rKGWo6tyzaIKMwVwpGY3kazYFglS6t1KtMzutn5gtRWqX9NoRbp/bDppoAqUtzsln8sGXWDI
wdA/Ii8Xh0D9XM+66EfaZz4Zsc6TW+2zmuyfgNJKFCLdoLDtLGnn2T/9o2i6KP+4MpErie/waF00
lwcSKQEuMhPY63tJ5Zvs8mGNtN7tulTlbX3YLYQG0tNimwRDjCS7NlXGwOzzEehNm7sd/n+KTykX
ozj8QOZpNuapLQl/RYe9cuHjf2GyZVOVytBpwUl565YNghRBZv5Ah5EwkvP9lYaa/jZWFZVMbyXQ
2CucsmhdIm+B8DxYfkwOC0MrW5tQdikJLrdNXwBsxSP50mg1vnhS4Q8k8MnjfEgqlHKENO3PlVc+
Qo33arEYg+61lW1/zmrzAEEKVs1hIXsDs8T6SNQJb/x1ixjE5655npGw1Q2dNA3+SZWewc0d8MmT
TKVYQDlmx+bXV8hCzPrNRdVJBKDEVda+k1ga+6X5qZORrJ5oCFfGmX4oZar0yJ28FsGxpFe6L4XP
M4ZmDSzvSBMuLi2Mz1b7S8mCAGsVnzm5rmTSO/aX8EgVZpE98+zsJ/q9YMhMGYiu7JVXJLnmav62
97qUck3CvNruGDN7M5T2014BBI9ofpPau7nyN56IPeF+siWFPcFkvXOwBPT9tgSF6Df/CTt4CCu/
u0Q+aytcAMIfxeHt3aQuk8W2Ky2+ZRU3MO/8HKAhruWz/qCNU/e9MLKDTIC664lJ/hyoibOVFHoC
frbuKd4irWi/3YfRfJn33w64CsAff+ZvaTHdb4NJ5gBd0JkUsDSB1CkwIOpAV9h5Jy4xGJizv4NG
ciTuXahYhtjfI16TZDulfYZSc7U09TXZGt09vXjFrGi6Uaav3EQyxP3ueu5n2dspTXVBgMrjx5MY
0EGnFOR3I0zzA13XhCFxA5uhgycGzo40TjKHuhKqfg3I0LFYM1F7nxv2Yx/r8H4/Z3H51urQz4xy
gMuFBcoTgPt1hEauWIc3VsVz+0825k7DQH37pIjDeSwHeYeeIc9UOMajDgv7JuFTdyx5BF1QdD8R
hSqWjkP4jTuUpWV4qHohKOxSvMT1W7IN+4QfaHcyatXCmEnuNde0vGSlt+2vuTI2vLuDO/xbi07b
zCBH9WGuuXsEW08JRQkNvvuyopD+8MkjbzXBHNPvLUYtzFMv+nV1WQaQI3W+Z1IR6/ThAoMJUeSV
SLz9q2e+DRv0kGh7etF25UYAGENWFhRBR4VeuzVw7gwMziWKeelVzeYP/0B17g2zVfXCv+JzcTa0
KN4EUvLKratZoHekA+JOwb2rqLInjGN+CPge8u9Gp9b/0yN9rSgTRRIczIz8nzPNCrTAmE/JqMgQ
xLUqqBeArqMoan6uajDOmRWyaECxaaiSKIxDhzFEWEM4kHMsJn5T1ASNbhztWQWndApp75YiLSUr
jHjME4+hCRowBDBvEsVuPNOra3yGZgnUe9fJitDcnkw1IZcTQ8wl37So6r/f4BoUaS7MXDRfjmTT
3wSODQ+PkxP+XW6fTU7wUq2Ky3cxJmx46OLeWQycvp8fAcT2+JkOJnBWjKA1UPSphU4BupMgHlqs
c0li5dZbyOZiqOjXxuilvHhxabNv9pg6pbKcjdSooZDxn4k7ROcal0fOg21hDrMDZHH5dbTF8gYj
QCJtVMQOx6Ykk5e/nYAHrgW8+XljcJ3IQd1r69reWdePfMAgAz6cOYlOfgNfN42g/E63T2to5k+b
mQNPbG1WYD3WOV0zRboRuoajEGOFykEZcdCVocPoeY+3DJiwLFc02oPbGLiHrRdM13LVLYRL9LWk
9oetf9osItq0ZALV0VOCbLlbKyiO1zynPPhhMNdSdsWwp5Ji7d5Mqpkyrez+qG5Pr72f4bcLKX9m
tFw+W3LgL5Dlatrng7oVENmVupE/y/Br2VZuTPw5iljjm4bQtEXhU3dw0ADbv8EtV8Ly+o9OmGaK
ScJgY11xUhxerNh48j63cFiDb6SWNUt7v5M1/lOkurUv7vJIOJb38+zOq8zK8drW/G6U0CvHGrns
+tGioNcRIf6GlGgrBlzHBi4bVeIqg3J9IzywJ1hmLBJSBpstXsKuOH6k4C0fGL2cbDotAGSzmjrk
vgWOvJNGLf3AGDg/36reFWm8J95W5cJhi80VVA+c8oX155Xe++sQJFs7TwY163hv4H4l/UafKxr5
WwRn9fdRFrKGRWZlbipOna2vURX5RsAtzWQcAiBA3ycRj1PatDJxG5woWWvvBvtn9SNBVBoR/N7G
0PFvWzKp1kFC/RzXwQ7qt4zfNUFIHWhtbmCWgouNKAdoFb2lnwLXegRPulRo4UCVgoXTvBGPWK4z
8QPLGW5i6YVoUTiwIfsmosvm5WP6goNZfsfiyTn0ddq7uegsWayVkxTitu1A7MvIrXTf11rE5iC2
otay+Y2upOpU/HV6oX/nM6lp1coTKa8ShWE58h5ZMacB/WUu3ftH6K2kBiXmbtxmRYuU4HoI1QvA
MTSDCWpjMTW2Sr3iG5DEqJgoc2AieLHLgxAao+FGeo0nxvr2IYEwx3DuEsn+olpRNurmoOXEqG6U
7/h0P3WzXrzRIsdnVVP7ANoKLGGLnLlYrfows0Sy8euKSooPEXroEXQV4FT42YjdazWKeWbGp9bl
EsMlkvn8D+FjzJ9TRPkQm+QM92Ry+X2906llq81tgnmEmCdW1EV56l/kQMd6lWjoTyBd2OA6w1x3
8/B3dThpvsLdpY1IBL/649ifvncUvfg/xg4Ko6OLSBR8qQ7n7DbFCWg1OiV+defWf7b4xvSKwfaC
bF6z8Rx5Sf/PRhYZOA9BCYEzD7Qln50TPld7oFPVuXoLdhXt5Vid78WC9z3IDqLiYZSrE3ABPA7c
PcStq8xn/vGxbF1Jp4VqmDtZf1mBnZjr+Q/3Sstll28tQQUbN5LMkmXsZHY43MdHWI9UuuypTkQK
EwAi0kDb/1SxcvvJ5RYIdE6Y8nKcR+lHPl+Y3/Vfwc7mSHF7vh0x8TNfO7tvlK/IZ43FOdRIXvgZ
kSAlhvpiukECmspIv5apk65CkUZUUtsmU4rratm7oobszvBkNR5oCgdQtBEppoDe7EAHLAC+7s9D
52nQMWUrSImYK86f+PR4uMhtIYpuueXDrS06WQTH1buRd9T7udGQTarVnQyFk8VUu4CcWtgkHqw4
/hrNm1wIRsQKcyU+Zy7uRl0G9sRVK0QO4L7LW4/5dXi5E4qq8e3rzDxMcTyED5hf+ExqbpazdgBP
QjLaUpjWiwimzeuDgLrcOsWQVfIZ28j5QiRl7iuEwGuxUVy97fJkja9Mg68yBHdcnjUyHE0z80kS
5Hngr/SrdKJrXQonLKJ9bcZV8bXD60NTd5DdUa2XmbI6EWU0fe7NuyUg9BJlNseN1j07kAi5GeO2
urX9cbHEymgorwNA8WYDtGttis17jF+u6qtBBTXyKFgkyCeGd/A5ZiOorF4Wd6LQHGTE2+hVMlHx
1xATf5Oh9IcD61qwtVK8mZ7F2yFRYly6Q7hjcvmypKVB/mwK9VmavC65EQ8uznMRnWOueAFTHYCi
/OxkTNfiXxb0IJ5idFUw7DxNFl5+gA8RCbfZzPc6xNs+RDb4khBrj/FoVpHJrSwv8eYCcH6fAvvy
IDvdKWI5+qkIQ4cJdtQCInL8PGsiD1cZF0c+jARHtTD/nLabk2/Dtx0E3PiLKJ2r8IfUponZFyC1
TugIyLFuPR9ouX2Eswjtth6M8BEVrnxS+4zRtaBcKfcsrajLZc84pVUBkCjA2/mHQPsianMOfw3U
0PZ+tYaMBVy30eiIXzPjsCfX7+vFVe96uBsN+x9pVHgP/vhzbd167R7wXnStu/sb2iPvK3WH8wxT
nlAdUdmpsirfk7wmtxP4a5DwCra54ZutA7uypGmKRC+cAH+O+c4wb3oL0qUAXT/KmcXHew9DYaRT
Z4QHST0J1H4lbXXl0ENEMLAzGzDPh7S76ew/buCFHLtVtIyWejNnsysws5Ye+e3REnr1XJZqwxBf
11fBqGRJnOal5WXMv8vqECAXlISNEFlVtzJNAId7i2Wx17v569lqxaEzo8Eu1rIRDEpZkoobZ2I2
VkZl24DaDOasx6SroRzTVdb+whO5sbuXB6zcu22SXKwd2NhmdTlskKrU5reyIVzeHSukF0VIiQDy
R0b03Y3C08iogE2rTYmA/j81X1SaFfwc3UWWKnKA9ZczS8kNk8qNBn0CSIQFTToNMc6jG4zrezUr
zh2P7HPUQgz8Ybjou0BisbAxZdW0NgOHQRVcyTdM1nK2aTK5jSvR/fLcCgosdijTTihOWLucg1Qy
9nEYA7cfIBeoCGGb8HS1PU20R1Wnrwn2g35wDHMis2m3Fezbp80KLcZxhos9ZKmLdV7MylNubHmv
yu1moc/VxuIE72AFV9tSNtxCVl5/b/kjxvlZavk3S7S5+1TMalKNmR+um6VnXGyg4wCYTmV1Grhg
rdQvNf9YJJgyAyX4dxzvuPfh6fm65BjAOJSGCEXMZWYGEocMCB93W1Hj0c/NSrEDNtWocpE1j4DH
GZOOrMswKWBiuMr705pY0kB+QmIKe4u6908Io9SO7CyPvjHXTfMj5RREqqSWvr8/7N3w04xGiBiz
c50aDzMlLy6aiEppqMfi4hpWevO3IPi96TR5wRvourG1O/GwQ2eP27fiDTsaXxNyeXW0DTqEcAqr
NzSm29yrfWR3c3K6YTaoameMHSlWwK1EihS6eg+xggms+F7voeN8RGCvOxc1R7H+K0AVIovJy7Fc
Oyfy6WQU5hsft35pfbunZJDA7D4/18KOnLx9AI0txPUo+tgf4bUNZeHwqnx3PFbgp+SbFnsAShn3
q96H84AOpdSExNfDmU41HeD2YZLqA9NT2b4Pqp50wmGzM9611MA7D79Bwdv3za/ZkGZSsJoPrJyU
6r6OaC3t4g9yt5wr3g7ahmFdA5juYohwTRVqYuaoXIk2PKHKjgIEu1uQwORflMt9WzgiMTejSeAd
q/kYjQh0it527FlUxjqqQknbg9O/afrgrDcy4lC6Drr8MnFEd90PXkdtbCUtzsM2uCKnXCJI255x
fXvVfF9pPgltVKWpQD9eeHxko90xLOv/cLP5j5VjHhOINVydPBTwohqkwvJGPVsyKJmTt+if5oiS
/twpM6gtCO9vjKR5zW2J2ftZZMWkJENenowYUlZv6eYRWbMsGQHQjBTY/D5RoyqE0QHRFyV0QYT9
ZoRrgjkSCim89wLMw2LTRRl6rLHmTd0TEOyImFlbvIeg3e4TelvjUQX2KkseyABfQAc5ijHLty/b
rVesZv8HQ5PkadnwUOs7DqIYdpkX9yCSYkk1ru7s/QsxpqnvPBkNkV0+RXcCzhEooLoGGaNIvU4s
ucFZav9cLygO5XaJukilvNP16ODqfLG8PaP/6OqX9w8EI80xGQoa0hKwpCU1oDT3hCfo7E9XMQbS
2l59/xgOvO60L2EX8jtuW961PTN2x4DzR5bv8uJiIZ9BWRWH59J14elH7RtFbKd6ARwsTpvLsFs2
gWcRFOZYSEIdQ7Sc+sHjlpWSU2PiuLrFZVjtgsloDoThoeQbyF2Y28Uq2CHFgyJFYfjYyimemB1d
2LD0wMbeSozJjzCUcnP80HjEpvodeQwmVuVO6j5+j7cRnGYbQ5jqyP8pHXwXq95cMEF4vIvjgmaE
6iclfmGuFjuS5Vv6ax1t4/ahlcdOlNdbK607ArLuCGlTsiZk0BKg9BoudbBH+whlc53HBNLrqdYR
zAGtBQSkg3sdUy6MXLFKYS/RQ12GWBg+CR+prFeWx3+WZ0+8SzFNuDzFo26IpsQXndgN8yynLJdf
RhoN3WGbx7w7EcaC+7crSsskO+2tF+jzGdd85rMAxT47zMlrFGw90OUh+dIrUrgLkbYA0KY+mv9s
m8OX3RTnPWC7mnH1i1rEF8jUEA4FHz73oq9yb8+R0Ga7nqcp0LkwaIwhClN+ef+hghQ70k/Y6skO
L6wT8sWm4JCZdJ1a8lPF4LiPg+FJk1IcUE9MzEzaWn65vhC+hvhYXa+19n18+Xv2JpLZCi4BI1iT
tUVtV9BlwTVgqWU7a0Folz6D0gribg7GiEwiLujPKHOHlriXICqzmwwFRK4QIPlL9Kur3YZaDAtP
F+BRqwlrbVbEt4L6YSzrw6a0PDFDjmlb+3EJOFaIArPoPgB+5hhFkDNIWjleWKSd8e+Ic63nURLv
obJnMifxl7/v6SlDyJaaMHh0KuChmKgCqTaWWMGWe4vYdgMiNinOnD070JsoxmmT1j6h10AoJiqP
iWoAQIFU7bjLGpQUwNaFLoBTSEnl7xGgJHCfJZlc8YGxc1Vo3sUCyQzFFaBFqy81PLnuf17c6A8Y
R227kvyMbne0C6vVmEAeJdj9lk5OVPMuNdKlR2xAUnpv/wFTOlckTQAPezgxpoGjfzxyWSlMsSew
aRUHzYksYKjX+pP89mr8sY9RjIxOCPv+46Qrx5S4FNjQLUqlZdq/wNBA3hRQPDtGOFDk3qNNVOi7
cGVJJTWKRkVX/j5F6q/1HicsZvi23/SL1tXHeQKmgClfqz2kK7K35zcLgShptx+NQJWhT91e+LRH
nIKvBzQjFirPfLq/vKfUlS0uM0Dt9zC3lQEGlxuDNyIKsX5UEad/7CKGTEjbVlcgYM6n4U0wpSLq
a+wo39UTx9m+wxTv1IpvXdoCKTGYj2XT4N5NgyPzjxdprLGYS8KN/JhrXWud+cQLUm0XiZY21h+U
k3a1TFBY6AHmTi/ToA7Q61iJJiQGfdsjKcPUBEWlSebYnE5iw9X3a1/flueqp7ioNOKQRByT0Mhi
BvYKizC6yYFV5K5WPIO1uDBNgkw9oadGMZs3uvb7MW11V0jkXGZ7rCNTETya1jWP1vzNTKoJ/KEw
QEHpNhV7RX2q5RQS/is08KJaayhBSqlK84j4q0Cq0nzAy4Ji1sGpVPrAvK3JEM5SwC9MExu7j+UD
yNPyK59qsJDalLGG2Xbt1OHiKnSwMETdoaW3fsYL2pVAwX7T/1PcxCPSH4XCxNpBYoFnSM8gJu5R
lapt/frTSJV+YEKTkd7jgVTkjhZyT2iRyBvTk1xKo1GxA2VQBZW5sJ1+KB+M+HUVVtX1AHC8bSPW
FXKCZdeQjjS8KhoXDWRfd+Dr/Twaph47b3u4qSW0SbGPdNNqmBIKDtcihgZb9Oo5Ft3Ge05MLeIf
k1NsQ68Apd1sSqAWXGN/ZNF7QQP3l7JL26n5nvYkIFCgPD4Lq0Ow04IqcjiqxtHbIkMkaDbRIoHy
EOLzz/r6u+iU7oYJFX27HOQnxRq5sNBNqxg4+23ISVO5gVfXDdFOpcm0T4Cj4G5y8FXwbDtFB3Ir
gF/icSEmF/0K8bG9g9I9cNR0zBfkI9RTU0VQDrF4X5nBs1ASz9hsvG8ZOslrvgrui2/Jqw192lHx
3bt1L0ZES77hGqY+cdTVLpTeNouO4cZyObx95er864mye3M1dGuctap4nnXLFaxvAD2Ppy/gQhyr
Z0CpejZAnBe1M1Jp+CGFS5I7bmbutdM5h5S0j20Cx1bTs2tXrlOfSL2AsTlGzxc5Brd5wtN4Jw1r
VpjqA3Mzv9CGxbzPq/6dyI/9pqpektP1FcO75lVKo9veP0NjZMX9g/AhgOfdzidlEHuxgRpLMk7V
P56dTIaXdKf3qhUx5pUm6lO+rzAyg0ihNbOaVKDRw8KdDsoY56f6HD6iCEHQguNqm2E0ZtcQcXZo
RFkrbvOzvHR+MA6bwUNfP4QbdVKDDf1sVjA/ts9+7iw4SuOFRyHXjN8NBz3vlEc1PuKKZLP2sT9N
yMmaoGfSDMF/L2X5BRNUg/KaVwUXxenbDDtu8XpsLCkZbOze4tqF1G1ogu+TaX4iIOWZqDuJOC0C
t1wCAwee5eAu+EEec6eLFuSW+i5/H6NuzkSy22VWIe+3bxL5iffkYZ0JAnb5Kn8oGpFOADAPwEFP
X9EgQO76LqhiqF5E12x/1sBdTW7Wx6uTJFc5UIAY+BswiC7Lzlxu2tZ7orEZdZwni6CjltfkQVUc
5jsZrwTkLK4RexfOZojAf5JA1tK+Tk84+2iubvtUSdsNeunG/ZKm0RONhRViCcIHBeUKhW4sZLp1
YHWOzE372F3Yare+3clzVItRjNPbnkSCdvmIsUqecx5kaDlIKfqTG5R35OGA7GeM9QcjuOKPp1Rb
EjdaRsAxZe77oykFZOTAVb8IM8v8PlxH970ROTptpWRYPFC0bssSpZSJXI+8ScpUnjNl60vTu1nb
IdaiwMvfkDJWJq6bp+DJfAvKL/y9VmqWfUBcGQJXinBDLHfl9w4raWIFFETzaRrehXpe0miiKAWA
oBhmRgXb1CmX4G8QI0j3Af9RlSrjEl/bYI9PAfAz3sOvl4XoZw6AtTQZjrCND65bfm5RAOTUw0Dw
UlQM7Ckfv0zUCRVpQr2NsPKU0oA6UtefnAxtgUwETM/VWxcAQYYR6kSBfeptZkmybXXM1p2KuF/W
q10deDyzIej3CvDJQ0tgWsMZ2cyJWFcY3Whbxbb0bYeqsgJjp4PiEBAuB6AgHT2tbfwor9O1Gsls
MTsiTHkRzFzLK7dzzKTwko9U0e68FjJGEwb4UFTs+mQp0nSnkG7QqkZvFq808b2CKeAuDJzfN+zP
XXDmS6/0MkAGAXtWKZEoGI26VPDHsPFOUEPPBDx6IN1xD+L0sk8X0zpiOle2Mn0OJ02W/RV2UIIo
b9cPuBUxaLAyqLsitVxDfq4TLk3XE8BKmAHSYApGTRuXuUrAR2cebMxTdtPscK3WIhYSi/8pzLQz
H/0QPyoqu6+BLEZIFCFqfnnETshw8ya9vX61Y5OLB+vY7dyVD/ExD/3nJt4TXaN20obue/gdRWqX
vx/J1bb2GNgD5rLgEIGq0Jccb//43hSFCgzq/ql0VF3Ou/X1HCVHsLJIQ+oR9tKOlOF0YMkGOc5E
A4d2Bh18AVq2AiEODBxH2ent5RokJhfE7EsxU1x+Pjr0L7X40hYOPEgtYQc+64pMIY7iV+fgzdRf
OQzajZjtXyBl2/o+GaNCmnf+5L+0FuvuShJLk9zVbAl9VOHdCCYG6IdBNixhl5hJwBIzlKE5S0jT
FO+w6tAuVyu3mYXnknMZ6WeX8tVKOmgDE5Oz5/KhH6eFwgSxvvNXDUUUyulZT1nvWz7gayPx8w0v
Va9RHKYOlBaOLyVE6GW7qAAxfnD17PEIbGIyl07BHvoTyKZUJuETQWBQHTcnDg4r16ovTGWOCImy
D6iP+EDreIi34z8SgaRT/ZGtar6yuJx/tGiHPHfEqwKFNW6fT8HcUMorAH4pZ8/wKFChb7oXzAZ5
Ybnkmc+38HYi1NJ7ng2ucBJOWTmUBjZdRJRbDDAVa761ej1mJko0NEhnHYP/lV9YfHHnvABcNA2N
FMYv2ucJPVrwyFkk4EC0BbwpsP2BdGn+8JccQN1Wc797cKW/4/hZBFHMSJCZrpKzudt0eHgdMM6A
rCI1xG1vCF/o2XtC2ZASpZo9ky+RbwKGJBJtaAPolcsSZmcflzx5aCoXdpsvpEaFauV5MTi7jlyA
eqhtLubeOhkMR29hnqW+Y2eFh4/5eH0WZjWHL6Jvs7G5YVouNHo0MB5YdtzwATfDQ0zbqruHfgiE
YBXPwdWmbRvrouXDI9iEWlTlvUKxwUsMu/caureauJxeE78JtLnEsCrEw84xumlh+7sZj248Nltm
btg01GARLtEQzGRBedsHitb/MU6X8JkL9HwnXWAyuwdmrJn+yBa1ARhXZb9wjNeu7GSVtbm5h7uT
i+GWmOc8/C0yPe3+5W1OBruh8ZN9m/eCMe5lnr6F5ufdidQrPXmllDYGk9GDYU2Tnsz1xtya07C0
+4ujHJ6rCVWtIuJRgosnnKEfVkOWVMixRUK0O9EsNzj9dq2OvI1AcAvIrJIzOjGcb4TjQAnGLwro
iWYjEeFRa2dE8mxU50BO4HPp0a36K7Xao2vM19wt5ZlOQXwJ2Xrda3QLTW1AvhPHnBgjqNfSDWBL
vOgExaZ8Z9JC3LQq58Q/HEV1hjSOuX/Zco81BVmG3wZBHn2yi1Gv1SygeNr//nclqL80AcaOEW1/
hKC01gcO3mzad5I5mhhkYzhk7nBtEMzKhU6SJBUxsEG9qoKNBel+65+MiXPLxwv0OZnAwQ5IETRj
8NX89v8+KdN1z+2j9hc0IXXwCBVyTpNTO3zYjAY6IbD9rnHqOdP+knBdM2zx6PPyaTwBiXSPpTYf
NmZvYtTfnSxHWLOv5IigZ7nJSxmB7CaG+Jx5I9y/snOEoF9CVde44fj31iBSWlNYraLU5bgm2xjG
d1cLLBAH+bNDSIW9FEJDiU67CX3TmD5ea6PADYBmfHccWmVJnZxw7Myk3HG6/JusYo1/9pXQhjC/
bIrB6XfyR3/LhIt4dse9wVEPURuuMJ+tmLF3L49W/uLaZva6EmYwdHfknACQVogHpXdskwpuH9fu
Fh318wOiacqErGMmzBM9Et2RXrKZgyQWGs6QB3UsQVssQonOC+21z7n/1DpelNpuBsEkg5k1sN6o
6Q8lKglSrV7TSkZJONIdHa2zQmZnl9g7nLw8CHDhHQ6p48miUUrPIEy7vwVNzdGkz7B+MoCfi1vq
x9LkgLIrBIBVH9V6/0B6MMp9j7gZ08zQERYiWsh22nlxVDKxiGdZgSLwSCdZT1/dlhpMP23cbxtz
8Nr+Eu7KWwU6ZSP/EA+rosyFZqUjqYZj0S3tULvBL+qJSEmNfJs2c9q5qYJYP3s23ArbX3j5l+HU
PuqSLPuvd6BMumFvDnDRmwODB3ou3zbdnLsQsq80N0bIX0FGpJCdx/bAMVtdPwZlrRLt4NgriLZv
bQb+XcbB9k917iEkvXqRrYj80WznNcjcw/4DWIhA+sEw55EBI+6cFcJf3CVoLwrlTrOvjTDLagDn
WwMxqaJsU0oC+XPw+6veGmliiWror26hLkyUmZoXXg/FEi+YGMYh//H4etEpPd3Gl3OWbRIuI+Nz
Mp/Kv1d8zg4LQ/Qn4W3jch6988w/0cY/Ybw6yEnWpTHsqi16xxIz1vZ276R4mSLkj+8aSlH2i+lj
/w5E2uqEa9zQsVh2htIi23Rp1YxOoxqIDEDRBTn5me+ItQ1sR9lljIP6JV5accWGKI+TyBQZeMsz
IF7N/3IGGStIvGOK8eqnWNxB9oo70PqSwiFjD71R1pXYaiPkKYEz6MNYjDEsuD9Hdh70wjtXB8mg
9XOOAcgbezbmwpqEePgKuoAoIzWdtapRDgNwiRRKPM+7NIYyeLDa2yhPtPn39OE8gz+K+Bs+5LX4
s/N9e2GCWuMGb+jU224681nukA6aOvNKMnRYR2s7WXaTC9IoPQyJsw0Af0poYnt3sbqacYr1e83+
Q+3j7Gz4C6fxwGGfp7u3n2VcBa6rVAPgfajvNMP0zQKhAX0zGqnetYtrMxJRm+cfvoEA8CzGYao7
iRxqbHdxLpffgclaUlAPm7khnMHuSYGilmE/0iM+znUGnJpwxZiqe4ZuW3DdcIYktMqc44wOJ2u5
ceYF2iBXFK9RWSJB8wTROcHHpkaZ4BifANV92sGxcRICe1o7OOMAblhGzskBNWdWLzVVPu8KMlgX
dt3Otb7XjN4uL+7xKv35l0QQxsdq8eKVGUc2PfhycyHOBwkh7pXwQySGfxCEkd6rb0ueh45EbhLR
MBl3c/dTIqHInYo4nLjvChPRulSuka83G82RmdBs+T+OOmgPVe9pQe0JsjtGYr3fCl2iCKjFRhyL
L4Gof7Marv+RM6sn3KFCnj491ns4xHSTXWoSIGq/uhB1tZffwrWI8TxkJ2SmSGgzbc1ZgC5Q4r9a
F/tGHBQft0M2bXEHHmVHHFYVswTQ+C72TS5is6JBjFyIOnpmo7nXUZ3Uuu1tg6KFkB5J90DHLqM3
0mGO2zrRnK287Bwc/KHkXYWjFxa63Gfd2gKv5os3VjPccN7heMwQNr5wa6z8IxNoIhXlNMXjzt5P
2EEDLPWF7MMPsvrLAcILIGpaPmfBRwT/6Uf0xfVQOs/NfnZ54G2LDEn4pXqm9EUoi9/qSG1esxJh
1R5BRPOz9zPycZJ0+YPO1BFJ44d+TT47Iu5TIshwkVkExw8Wcipa6ptjBPLaW+pGNND3nerfpOAc
GjxLps1IOx5YzH/xIxD3nTi7ArpUBS5qRfzbozAK3VdcaRc+47cTw88vKhkdefbOHW11wHpdcIGR
21m2N3f4+z/vWzHDnCB5RuOjCtoCqf3ygpF9k+BlgWEyDKl6DzrS6nygpDNKA2GL74NdnJTbI/rh
JMKsmXSVWBp2Gt5yVZP3EDs9mPkNwFT29frbkEI6S7alZ8kIAAf08csyz7Cx9yzDGYFhyCXIdwiL
7vYjDctOrjoKkB9g2ENO38smhASMMM4R2ba4mSgCBCJFFqv7PCcWXhAlsLsOl/CdZkCEFiGjW7mx
DhPsbm6BnV6dag9p26Tx3kzDKP9OD4k/WZS2VENaYJg/BLjyNp1ksHLWBgJitcx6C+7zK+c6XRpG
Ex8RpzAEmbJNxz469nJFjlOxS9GffPp8+/jm4ZxsQjU9q9ML9JcqNbNRieVQQ8hvAKQEpoBiydSH
IES0KcYQxdKKveYzM55IyUUb1H2uRfaYjiEGKhzkzEHV77vRFvzFjCn3ftXdfWIM0ynLlyooih0w
cb7WZp2HUZaV/2imIyqZq2z5DwDdXKaU8Sx+F78omgYLne8um6AHqPtM1VQZWdKQr4DATl75hWUz
A48VOsebKb2rnyDFSvfYPqN64xdB4Ukw7WZBsx8/yu5EFm4G8Igf2U2cz/AgvKSmwj8W62XC2pBc
2/UEqgKSFXPRaU/BMrCYOW1Xb4eZUg5fZdjSLzw/FDPS05bJF4h7GaKb+1jd1yYrYTJs+sXfx07Z
zLykZnXqXxRECNbZgV9gd1pPjoZyQAbMWlR172H18D7/ShDsNfAN8qUKzr5U7dyTXs9pKl+ZMIlc
fV7isqaoFryJuEgzZFoSCmBXOVm4TTdTSf7fcEepDITdPFrllcGyMf/28pBXt6kfD0T9eXHd3E7O
qo3mp2FuyI41IfwANSs1HE3Prza0mYYK+QrH0NIMd8Q7ANg0DNrQk3Pu+YT6WxyUBxTa5ipnZ5iw
E8hWB+gMJI0CRqAXDC8Wh3tBWu5UkOsoBYBQcrmtxYxXH15cMhYrVezFjU7OlbEtAMcjqTZim3jB
JUI59HoLFY5HnMIAJtLf/MxCL3LYh1mYPxEaPyPM0jMGDXSPpXU0FFZEorCohD+zjxjndw+gBEec
/lKLfeB4xY1jDWJDAv+uh9IhDU8SqfMUsycqyq88XoQ0+PZV5I8HHEROvht0dNQDzSRmGgXqVqQy
v3tFVw3AEvjputATgKQmjbxqGOK3QirzNuTb26iR1SYwC/CaAfPLRYjZkE2lv8+ly8XDuRsEbj0u
/QUIaSkynM7DrCC7QXP3D47hx8ldv+5bNhn8qffSEvuTa0YGd2bihiqbbaRmQDmWVmvIUc06MOML
fO9GGKB16F/VHYARmKP0yNkAuYRThFf3H9D0kZqhwWR8VLzuBjNHEC4oItMySyiTbqRl2FR28aL4
M92n6mfQYBTTw+j7agzEcbpcg01bp3F7DBsNOJag7yN+akFd9nlLxreten55SbWSIpYrJPOE7Knd
qXXJSA5qcLbD53V5h1ds2+1PDwl0TQ3PW+NJ+fVkEO+1ZYn16gwtH7omVz4tnAY40REcBIQ5WB0n
Yut8oF9zET6GD5FQHnYkIgMQ4HdsQ/3CHuc0EvN+4VLCVFiJtdXcisaLtsrIAMT0WLk8S0/8wSP/
4/kJMnKVpJalWEz5cUaDnT7XY4RWBHi4KcodSnNUYmpjeHaNRn79j+T0fSJRf293ppJqYLtBYHcj
/UkRSAkbTJ/xWweV+C6wPUYmu5teOkVnAXWxLe97u8ZlKC2CeWWHvWac2++WLx5MD+luxaJ1Dxtj
1fDgPNYswgsDrIBfGb+lPVHge9nQaZ7bzqsdq++4ehHGVie32GXJWMCEMu2V/JvvT7g28e/AO01t
M7Fw9DTdaSB+1C4eXw3NB4ozXq8wbpLdKvFxT3pDW6ASp4v7yd1K7pVZC6NC+rOD1AGWoDVvYX97
EWOSQ8XTBkbMVnPS4OOPDnYXpS8Tf96ifmFA3uxROT0WKKVHNqzekkz8+DK3ntcXvHz8Ptya2+UL
4ZW+N0Ot6Wr+tkvxwnqoH1w8rLAub8I2e5nax+19+sA8jxMxblGBt89nWik1XXlFk5zZLz5m8Cvs
b8lF25aLFnFHSbj55nD1aXItZfRQMmo6j5VAfJPqWY8dElfSHwbbRarqj0CFAgR6pWPJW90y/GD+
2AS39nK2syd9E7tJdMlE5lJYZ5bEyYWyMBW2cU0XxNY0yg3CCr2O9vkNT7Js37GOf8pg6MlOUWnr
KbJ8VlxRybY9+DrBUd57o2yr1mDBMvyQPZFYj2ESZkzKny1XvfimNx3HhLEAlGqDSU4mv8F0gM38
KkRcUNGwxtqOmaEb5MXnUyOCD7PD6iGhNeVqfhNJD255ozOyzqdLRTle/70VxX1jH1BzIRv6fUpk
NUFbr4Ou+WdC9s8mk+/KrJxQvqdBsI4big/xKV6/YB+oNuBX5kTL2Byv12dr/hWq1wUtAklvwHPa
50SZOTc0L/6AO/F2SwDNiw5Tl1WM+vdFktcrkB9m6+VEakYJx/Wwf/yW2HHHThikd0tg/ioF9aAa
MVEeha/9E+W/KRVtp942BgBjsZxY1HJ5heUgIPNI0fjPuc7Jup3auEHgokuxYklZdPSmrZ+h8moh
qP7UIej9WN2ITuzJmgzj/sQmZrj4cxY0qY8J8vxHGMFPzaQV4pHOY3RRJqxOXr9jWZshKSrcP7MW
PUq6BtXqWgH+Hq8e6O2hXaicgmdg6Nw7JZyzBa6Ogex6m9cNBW+CbyjlddY5d0+aIWtxhdipgsL/
JbTOk07Se4fgJIthB4iPci8EvVpeZH92nbdb6SIV0zEppJUAH2tiBu1a1h4zpIlBOdU0PYrM02d8
vmS/IGoFCLOLQbHrCfO5UcL6L74iNfYk4pO36W38mx0Fi278OuvJVfYjmGNU0oOTkDMf1T+/3yAa
NQ9OZksdYC19N4yj9HvFrXJDlueHFrpkWQbz5/8Lkb58m6OYA7xzbwbopoU2iPbKFA26mHGslmr2
2gWKUIRbqzjowETIv3pIwk8v8iwHN4934EV09WOzNDxakpUkuQwTs1oACRbbiqNpmRPjCWqyuySV
O7DtBgqmpyj/khrU2gePXStqIsfXgFM/rKjamvDrukr9PTXC6Tc0hseZQF1LleLvBuOfeOjeNdIa
8o++lAG23D4kc9fwHiPtmzyTZ8xHfBY5GFr0R+wAFFVyrl6wjFVJHjUw1vbDqGcztpJq2Q2p4Gkz
uapRFQ508ZlR/qh56P+sm0/5xaroW88Xv7mfl1Mye+7joBrvJxssWaJRkb5mu3LmJJhyrJC+FAzo
N8J82aD8Y88VlmNtUWig7K+JjcY5fatY3uUXRQWrrEzbmhZJEhmTk82JLhSegw68MtgvZxSp6P5l
JG6IE8x64lPY/mllTiY2Cs7aUQAMbnhg1w1AXm5WKXkBbWljxzj64btN3AO0BklqvuPcnadZ4aFh
yi93pxYGoVcXF/Fpp1ogkg7SgjTKx+WOAeIQpdWHHIGXLDRRi4ckkqKhC4J181hI/TgXOsjnaVMY
T1IJmOLpVqFgU5iZrPMgnGEL8/LSaggJcYDQH4BFs1vwB5iCXAOwLj5VxRQgwOIDoBtUIwRwFjAd
uTbmNpyAoOx5CjEDaur/2WXeAJptfuVxi02XQvPAlKsjftS/hOaX3BQHXom4QMtogMlwFJ5Wrq1T
d3VJDnzUYujNZhq9c/r93W2YHPSQoN/jKPJe75HUuXcpPC+bW8YpSbc72ul2AT+5bHLPxJhVK5N9
ZHVyttjORZHc5ZMsvnCVQu3kMOlSnwL+Niqd8crUKMeDQGqXOnL6Ra3obXr45+0Y0+iS8NsI2FmS
bK+lHRJ/lkjNUrNDXvtPtPzvIPK3QfSQUGOxbnMz0sJIuTGtNO3mP7075WdIc9zeeMxfQqWHR5gS
MP98lM/yegn6B+mGtDVWJWZUElI8hGB+3wu2WIJzV5/+0H1Zq6uM/WvvaxB0UEFVPHHAEfw1YHND
uXR/7LA2eO5hJ82tSRMaljV4B4WfYX8JD6cDOiZ6UcPwZ0tcbzOVr+0n9EdQQq+CuWoVcA8la2F6
gWoGAmArwJFZjqYQybFcgJ7dcRYAk10WcqMkNo/01ZUoSSNH13juTHUhz0CaVhs5dgXhTCBLc1lB
SE7W/TSwHhixuGmfXzuz1PMyKwPgdeXELuFfxkpQx57oGlfXhwbkFbFvjPkQVxatqbu7Juv3Jafq
3iV3JJhvPV9UK4inNxThp2rPNSVwhk5yDFaw0PULFc+X/LDdqqPFDSDTNjtoCbW7qhNrMGyYtvCe
7E8MXrHiEKgZisrHrXv7S0/XaLnzzPyJ6FUo+xd/nl2QX9uyi8e9MRn3e9/GzAHjD1BtizYVH3lQ
ajtJQpKSXfxuJenYivF+lCGckGQPfSJoYf2kEdj1jlAkV+gNIGm6ojTk5cUwEAPN82IXmbrAmewR
9Ga1Op1xctEQfee/CF6x2dTltB7uH9U4wtiz2fK8LxGzu6GJrx2iqdISy0DFXWi39dez5zUxv6mM
nXmYlMlev+zyMI5fpzkynstr/kI/uutf4rHADTMrap9dcq/pSO2H4afCeBI4fNCVHz9LmBzmzMT5
Vb5diqfGLaMcbIhG1G9mbGHXsz0Y7Wj9eSrvqV4HPMtqQZSzJdUACu/WxTgY3yy/kvE83RoIiC1M
34FCT+wO1rXftKecwFv6NDvl9Ox45CPH0UOqHQk5xNM+B0yybwkV4c6lvOc9VYxR5LEI3XFIaVmp
36qLAYPeaByxv7p1ljNr4dt7DGh0nWmaRbBFNj1C4ahkBlXonIiyWXqp7M/Mj733mJmReMcsuOiw
AI14TYzMAzTQQ6d4e21+wbEp104yiqxPoXtpCmrxRH2NNuoP4TKEvJzNhqeJnVQH3rIU8jlEnlnm
wXN6iG8kUO7FmgfOc2sa1qiW5x5qZpS9MQz575WgQpbWZt6tiFrnEq9BH6xPuDFiLJ+M1RVjySZY
vUj7bkP63fOmJiqBu3bffyF6aP7r1OcJPveJHs1YYT2pLKy35PUm8+w5tRDFelaSGrkOPX5kb2aV
cO6sKCKTlFXBrQjLm0ZmwEdxccSObAb43Q8NXdKKdBW6HSZuKyByFQ8Z82wbi3XLp4FExK0mOzKE
eT2XsjCuxn8sY6ehhyNvg6GYMPkUqUcvFHcjBwKK4vZ3+g4vsebCXg4rwL6zgnfLUat25g8+PD2J
RKvSXDxo5Z3sj2YomkAzni+aMms7JothOuNpKuPPVcuPcipRdD6k/67Er3AaN3XlxVreHrSW65b6
gMW4Uj/pF3I1WswxBYMeldPh0zBnJfXlgxxue8ZSLg257SpLqMw/+3Evu8bJLeOFmcHMh93hGadr
UT3CkdyFVAUy7Bmfq8PYxIcsft99Kj4w9uJs0nRUlxLgpBQ9wz/F0cG9s0vi1xm5jS0ZAhwUbeNv
O79u+36rh3Pf8f7GSCOpxbALskZ5jbbSyYyOJTpvpYR32U5GcmSzlMfXjmZuM1L7tvqNBWCYi/Ae
YmBReqbPVKIYzmjfi11/nttkYrB3kfzeHhIZ8MOG5Q2aYBC9vTND9za+2CYoy5rbZdqcLdcNO9L+
RJFfmXEY7Wmlg2F3wjQkR8VIbhf7Ht2CVVL3BWuL5LHf7obN7YQGK5NFCsrTHH2jfjdKBJtRlIBn
Sq9MdD2hTKXnaRS7rNJo/z8F0fLiAQHfw0Qj4dVm/4KgvJLpREskI+vQvecoETnJMe5azbG4KmjK
bMIg82Q4vYzWR+93eYTME0gHkzZOkTYWuM0tUsbVGiLpA88yyOXLisWiHhkp3FvZg2KOvM89hosU
NioMflAGPTDv9SMq2nPbnvJHNiZuPF21DX1Ezu5beElQvmPgfatHxdA9zIGxoTE1XKYJdyc8LK9Q
P2ag++57vp92EACYakTGt6H1FCUUAQet2eBAKYfp4HQVIMRlI6diS97VHel2giRh76+5tFZIa+5d
vkd8MiwWfMYV2wmH37M4280WvcqSHnV/QDccLGphuH9T2CV/wOHqgJaNGuH9oHsT1nH/bIuLLuDh
vH9GfYHzLbFO6zUL8oGdcRhHFCuWUjYuaHIvRi9ifYRSb75EkwOyapg28TZ3Ruale9on2d7EaPK+
OElY+2L94ZcEHPRMIxDMg50LZjO8ykqLWKq9ywW0ThHolEGUtu66Oa2tFUUGWPm/i37Gn/GBmCih
qCvKQmLROsDrMQqv6yVqQnXDL7P5havbmZ4J0xi+zTg93DXSMCl5uKH2pqCmFm8gtq2ioBGY8GCf
aeunoZTCREYPLJzeFGJKueePQfphS3lwphMlb5pkitwb5ghzUd/6rCQpNQPEOSD1qUCqeU7PBD+U
cub2SywPteJv+kEiI/Xl5v+SM6LOVsEgixmEkr7RN9Fe8/nkQQ7XKXv1b7aFKuA4BrK2SHO4XAcp
W8x0lONb7QVJY2zsdG1B3Nwao3QaG8mxeTmBAZkpBHQQfG/1wZ81r+tSsVilJzCBJHKZqJfhkM0A
x0mZlfRSZrcUZMMlxXAdOjKz8mFb39ZnE9h10Rw2f9Te+BL93zDSd9D4X95iCB3iev9Oo9L2S4Kx
HaMIIZ5uNOgKroBokzRRLL+L+727C5/M6b4CeDvG1vNY4GNB2sZdcNBXGfftby4GvSltEk6n9r92
9JFwZ4S3NW/TQi1sntin6d1Z1zetPRHZQciwr8YsLrZ4xb/9fRbdjOElUdSFJzbsyZKLciLi7OyK
5D8dDKpraeuF7H8/RKml47tDwTRKjrjYW07yMUhFNSVjd33S1GTLpfqm/qyFMOR8qILhYeVK/WOo
FLQ39RUnFXOD4wmOvj+uktSH5CFq4q5gjGYNZ7iqGpOMy4PjtndGvpGgkv/gGaN+AJNRmUFpEh1D
+//Xy2/dp677XSh21mgoI9iRS9H6qv2hSPJjG8VPoh6s7iLVA0oxk1Bedxlwj7R6SmfAs9vxOv0u
Q7ymD0zKi02h3fVvkx9lCZJYVKTLc053HW13avJ4e1h/4IaiEE9wuGxhqDOCxxfjsEb/wwrgeJhg
yYxeWjVWlXnsBY8WqqJlz6uDX9U+9q73YfU8VWHXGfNN4fNCHrA3VY8NXCdUyNkz6dXgAerZpzdU
mBBIF6wNYukOxIZw3yNYbvafraRoSer3YokeXkrEkrdP64ldzXApsRXgS8Hih2IAE+FoQmJ/1ys5
NhYGqvIxzyZ5Y7Vq5WuzqxinavTgnZikecWW1Fs3zxnHu1fLgdG0M0n1ylcxMtBDVOYPmNsuGIVg
P/c+zymcjYSIMe1TGrfkqlDrp8ZFwRSgvrWv5pAa47ypFJYL/HXNwZIR3Wp8iHuzoh+JG7Qf0tza
y86KnXYa+OHBbdiHU0q5nKwz5ZinNWdz0WVD7bmI+UBYaRbDHSxcgwWN3DxNFEbcH7+lX+3It3/E
5SFm12Kftr/Mb0zrhy55ArySh3Gm+xXRI+cn7T5vX12HBZ/uMfPcYeqJAkFcF+ocMOIViNYY94qE
4BTBp1B303kUjHZWF00lSPkir5N/84ZHaDFnU7fWOag3WSi12Tkps0L3PrQ4qEQU88d+w5O3Ttvn
AQTwz/+B2dC1Se/GxNfexayXbffBKaY5uwxcM4OeqlpYDJ1qwuzk+n6L27dHkCT6BCxLVG1Rr9Yf
RISbCfh11GoLTTNhc7R3QTrpKyJ5COYf84+WEkrs5tYgwhD5LVAMagxghepVAtdYQkyQXD3Kg4sB
tKF+BgKbmAXdLXVDdA/RDg8+Cmqpxlix7yx8JXLBbXOeeFy0Iuqktk8QE2nrFR8XXsU5+RE8cNk6
e6WuaDonvB+iWhTc6pj2cSy0maFQP3AnyqVgcvgB53ncskwz1MD2TVC0/IYDGYNRaxCgZPjT5YZQ
3k84FEyBRK5Bx7/lrhA+nOJJ/+P3oTrw7tJA5BOFRM4xm+/4V0mjuiv3JRfwNGEePzO0ubUAFT1t
A1NCErfv6OOKi5PWUcNk3QUmuQAVq5zNjC7UMW/MALEg+3d8wLvYifxJ7oeTob6eL+riCUFncdV4
x8pfZTQl7cR2HQnyokYF0vEhKcjoTZ2v7ius+Lzpvvp4/I/FBXJlXIXzAVVg7KMftpkS5wPGxRYd
dDDT1983Snaqr0B7PLeVBVt4Pdls4MZAlyYthtCeUs+l6Wj4RuUVTu8ku4DW3AVea/XmVvK1SlY3
bNtBHsjdodFRXLYvf8c7iyn47cYF2vQbE0qnrHXZHoK+tkijjx+1tpPPHx9mfmRlOvtymUUDBwGY
3VfXooIZTzeoArDEIWQBJIRPLCCJfADEmsEnNmMoitcVbTTRsqkwoMAB7bE+KJS1NGgMlCn4zSIl
z64CLzmdoe+AlXptDIW30Hja0Ter5M3x/Cfn8JzQSM8FeTvRAmi0iGPbv0eVzM+6Qxwqznr+VI3v
/ifj14KmbS9PB8EPbNACrmTjV7io9SJCIetQ0fnxfKN8PYmlHGPXNJM5uNPwZdzek6eeWD1gGaCM
f3Sy1n2JHVBN6vKxFi0VROGZuO8WAP5JJDQ3X736+NJ8y/tjjGTvdCXDHByP949HP9x3H/PLFJg0
8xqCq4uwT4yTg2n4zZguF6R185J2r5VMSuqVVXcImYGsJxd8Q/28jzXqTQ/CIZmAFO7YntTco8+e
OjyBioI8ysZwPv2/dyfycENyhlWszRnB6qwtCEf9SGIOeT7SwaLMM6vdjen3/bfYzBRbIeRj9+61
QqENss+m8+5YcUisaBEFGdPVko+lfMr1DQ/upmJ7NcWksUJ6XyWqyVUszkyhY/b4VZvKMloa8Wlh
EAYHEVMxIygYO9ehevmXYmJJiQK/6GHMJ2pwaZP4OeAUZX6GdhT/Hb3O0dOXYKa9kz3uo/v3C2s/
eJ9HDj3ppxPCTH9s/7R967olkY2MvBW9jT6S1KABnpQoE5UkntGPpypDhWIzcKHS9AaJsNbk5CLA
TYW2Utt8qipyWyOnjGm5wlHHLUaeMUHFJxiFPOXq6yUPB5Sx3YrBBfKKomeeleFE3SyzxGXy5SJA
sDt99XraAspfP9EoP/zFKGNJIJoP7+MRLNqpw1PiDcADjvmNHbZvO/Xrb/07RDoZoy/N9LmFHj1H
kF5EA2ykWMJD2w5+dRu7LJ8GF8NWlERWcNfYSbpVd6uT/b0qkCk+Da3nWVtZ3jBy13H5Iux+McHg
aM+CleabbH7X5JgOkooWpXduQlJEVXot18pjP5vcZ4KAcRjXoFrJD/09U90pv42mKmc1xD8eqvE3
kkLnJjTj4SS7LEn/2IsMozmYQXO5KwE2GpBc7DUDzwuJMtn71oucLOp5SlHVdJa7dHYJ7j/nuIiJ
d09GzchsCp0mxx9j9uLwZznH/7Isxi1yJ2Lw30S8glhq9XwGfhVhWNxwQKUF09uOGTW5SlKEDCCH
eKy5M8CB5lVWU5UjqSAXWWMgy2+0jZSAMRd8KSWmFN24qAglxi6nh5rOD3WIWfwF/Aa+OexqvzQc
arQsUa6/SNOoh4nqgULaMo1NffFIKSz7ri33OVrf1hLPTmYIcXtgEkabV0lmLOTFa/1ZZ/qW/QnC
Ejaumdayyonep732HnPuScSOphlTDF9Dy2vfwDfd+hZY+gSEBHCTXb0G1YY462LwUcjqsNzUXbMm
sPj5F9vEBDNkOjJSKC5JdKnqGHP4jTR/BWJDF1gOQkZAni4xCX0yUUWNGdQoJaqRVz3XWvBupNjP
TfNTWQ74LHvhes9ugAP7Sh8rWblOudzfxeWd6v+0YLh/Ndz53qldZqYX9V8HMdRjXuzGDHk7MWBz
b8aTSX2ROQ9CdsgK2SM/Cdf9UtgGsV6HK0vDb3uX77BZa7Veapzg6aaxH0c0KnWFvzBXLMm65zix
umHH+AIUskkn7QkRMNqgcvShcYRgXTVsSmODTrefFPQAl+JgQrVJW0OWQZUUb918zsGVeT26SFch
0WmhqvwjmKuYFM9tVN8ZSuEk31b+ZF8DpNPigR8jJZT+o+nnEzI5kHZx9ltPgBCgLDRUvkZIRz3A
gc52wuNDCqHMSzXBDn69BNEqDCgOrbIr8CHx1akG2aKAS4QpMXonPDypVUB7r3afiFmXBFJ6VA+o
xjrU8R9q3CiznDE/e8ERQa9aJSqoGV4R12JR1aNHZrXuXQl65+pq4Wt6quIl/63WqSA7ooq/bx0i
cM1eC9JtwFKKdklgbHQNGIDX5eG9ZqaY9/sZQsN5kksW4PW+kUQSEMI5xTBAOqr9YV08Nqjv7IsW
sCkiEyyH6nTG0e+UOx22Bmb3hsJjR3y6iElFkNVpxHWomostJpnHPiELdQ5GlJQDKazDj/5BjZX0
cEh+FlqnjH3nGyYGKhknvEo5u5V1GbhVZN/Jj8LaMzd0C0Hnc48b3plBLXrMmLrSVk76NE1pIT2Y
PT1+FQkm+D3fFbog88IxS0jcjAXcMWDdCdwK5ZQsyKZ+exJ6OwxQv2uq9uaiR7mgUqEOEPEQY+Bx
RNRMW2A4XVJoI/u4BpaFpwx1mKRU7FTanODq7nAFvTh03mmCOGMgR8X3/mGYWMHhJJcQa79A1P0M
pDiqOEWz5C9Zii3b5+MXpadmBFKOCPwRWyJvY5d2YZzl21KiHk2xZMNm6Yl6leSIbXD2baeI51d7
xe/l1oDHu9k6BXIOsWJkE0ZzzptM7swgWx6GrqNY8QMOriOwM63Ig0B9J7s+rt0WZaiQ1D5MizFe
OYuuKpHvohNqqJaAQGd1Aqpw9nLuBcE5hyYREuFese93QhvWoMsiiesmBOLwxFHru1x6Xwk/PVRh
CBRaSXiFFlSFvLZWf2DU9H99ry68YbsrT/zT0vcBIcFlgqwFX0hyNmLU+euacSx5JGPqk/YiPoQy
SOOq20sH3q/yUfuekOCuKwSIvVmHLJUzuCAlmc82Mm8sHjaHv32RdYIw21j1dTWTv7WN4aRdnbAR
u4+GxySndcNHB8xTZlCDjHBSPq9kZdZw+jP6DUjxSSb/03tWyNC/Ig0w2KHHLFeY2/EmTcaOY6oy
dIbGmej9fJiUvG7qzIy+jriZtvMl/4xm2qoLWJcdUowgWhEzV7fHyy+3jf5781L/1KzTdx+MusnZ
yOQa9DwPlzZTBNpPg2Pc51sm3Na0c0hAX1tWwBcTaiLySpM5GK2lPkT8X20iE0Cii2FICdpYbj9N
DORQU4qXDFwxZYlmDFbms5hmdEfaOL8DCqPFwAfqbGsxmeJlaIPBAOPBdEgExjIHTjW3w69rKZLN
dXUq1laJWQscfnmWIjBrqES3GN3TT/B5poPkc2DLj9r/1GMZDxzVmilXbInQEsfVfgU35oNOMwki
85YEL4XGijLlIm+4Jnj+To31E1qjU6BwwFzU2XCYjzzEyHMLTdUIuQRKrScckzuWN7DXpLXup9j/
dBP/YRDTAmh8RB0cMQDjopNu3p54PrK2tHZhuU1q2UwP0nuHIhJqvr5xZEd43EsMo0GnJ8rFQyV/
O1evQmjIXgn/YbwdadLMpDIqsZ377OIi5pLUBTFc3IR756NyZkLZe9a9+vZSCfjtfbcklAn7QZkf
Dw0Cs0QDiuGPQIDoKIXIklvnHb9um3WGgdQrWKwdzXPEuDEa+5DVr7sa8SF5w573H8VF2PugqEkS
nXw2xEqCvGu66v9gZsZY55IQkC9tI5kD8gL6bdXv0QAUBRT0GdAUzJ/sUxivu3X3Gaw+lNFMc7K3
wMRYV8fmyKOqWvn8i8PzrG9MErQVlxViDVDxSbAmpor1SoODBc3GcOFNNoTyMLL6P4guoNTOyajp
7BTZ4aqP0xECexOIFmhv4qr/H4WQD/MT1+v19l0EHLxcJ9skjmjTKb/5TzjUqn78QVQrwi029eyt
1P+914Ag041oTzByaUVJ55SwmBgnVBBM3+GUcoiWlSIQBISf8M5Q20nvdWu22uPrxl6MveQupTgg
4pXwPbWusGUePFVxNgzn42RqPj+fK5W9iGtuc7AevzunoHdwV1rFmSJCNQg2OWQhZY6M5OmV+/lq
LdySAKEFPp3YLiHpKSTMgl/3pUqvZYWZr+yJe6T1m+xPE+JKkVkmDHbVUQoM/wEVSuF8XA24kZAN
wK+s59JgELtxQgW0JoAfIbPKX4h/Y/TCheSBk377KsUskemS9kyOOsRMGvXjYEyQ+KPWgbRNd5UP
3EZXIgPm0Ww0AaufeqLu8UwJ9ieuwYVtYdrIK7rH+lB8pm7vTEc+sf4bAbnWKq3SGTvbU272kFEa
K0THap6VGuqakFBPDtp6YS319O/NsL8BGI/gqGlKEkUnxrvoFXFhwfhA2GaPzx/k1PVAmnomIZWm
R0lqC2i8rHAdxMJxYnSE4W+P1NvSHI9hul6TBm6KukZ2qS/zLX8kt8dJ7qXdnyQhsu8GtE6rQeKw
oxVjaE72Y5eXMOUXxwY3qExUcpGkV6a89wo3UZdCBXDe6Z5bvNWn7iMPJ/+chBo1hx7OX3yMGZlU
tv8biAiXY8qizRAd6Wn7wqAMaTKNhOlhiHQ0WmIvTclTAwdxdDuxuusFcys99hZ62p50L+chjc+W
UQSVXtGAY8G62RoRScg7S4pJSEzR9mYsMhmj+CCjeUhHRxkHTgx6rSIJvgoQ737LDtTKNW2ooLKB
V5qSyhkWZFMkt1yNxWtuWeYQIpTueHLARs5YjmCgumhPiYdFVFbZirVmwgJaba1n2CQZ4rRNWfWt
3bJfqRq00TVqXPjo/KCb/DuZDxONbrrHztSxMsLgKKkbgDycGCX9fkVZ6gTLb2qxZngPWHLQUcap
eZR0f4V+Eim3X9Mi5d3BEQZSQk+EKhf+sQzCA6mPmng8WzOa/vNt/ZIVeVr8/SN4SDRY3Z5hm00m
6qHHYLNuA2C0tBpXOrMDjF+Y8xQPQfxaTKQHvSmICjzF14Bn0AD0aji80532EvtfrCdRDlx3xY0V
/FoE8/57f9R0gc2SyjC+YYJ1MUrt3sf4RpZTARTnDQr2wMMq1PR+qdk7d5XXy2umxFV8Vu+mPdxc
OtXx/1g2n+FKSEdbQW4g8a0Ru865zPVXabkCW0rahYBhLcmXXShR+ini+a0vqIcw97waiXQ5W7Xa
23ey7mSf1uBD6r7fy9uonZrUmXshHpKLEn5vlAm/Tg1x65DmfWwZWl03wDooaCsZkUuasIgdF+oc
aNwirzd2FyThsjrOq1Ui9cWdsKNHiQY3ggUAazOnU06KhyV8J1e1dcsiFJVOmatYbIa5BVs4Dau2
c3AmuHEksrQnVMkwSW9ttEkoKeMslFA6bUGQXgrLEPBP4vFgS/NDW1TBz9vIi6jLcJqBxJpkcpPG
Dc0nrUFs9FLqPuUQxvIl8ifSKejJgcBzoQgKZ4RBgY2XzlkMfjv/fdxdhAFt1PgVrRy4axRUN9Jz
0PTR3ZYnJJXiwyEZpN2kMXU7snq7XBpW6UNYQDumeVCXgmLnj58HId1mArNuXjadT3pqjq6SUWcN
5nsYuLhvmSK2gRCVwqKZSCAt38MLKigV/VF6hgGFKgNH5jKojgIKJ4wRJp/9BOqcbXukFAHWdRvI
fnBUTkqRWco5yHKL+tm6Eir2IaPWliUmz2WEhzwkxH1oIMT+iSFIgOfCOWqWdr9HBVZVvzbNO6qb
scaq8J3J7DqVq0vOMJglF9UIOnJFLwwAUqO5MoqJ5NBf3+cgHkBaPZdWMjsP4eyL33zogVP2nkIj
OQgBqtBiGF38xcLKB2IkV5xrzBw1GqiN5DTO9gvGSB7tYT75g0Wz1Q8/bdLdNO5dp2A/wKgMZz1G
SqxXR/682ol7eaAPxXwxgHYydVWoXY5glYoTsJ6d3cWYE8AFptukGMbFgIe9T2P31WTrrdkI9zz7
M5P4pla7gTQYndz99Ymt8c7iVtXO+jjOHIuK6GUa2AB6KHSxwCMJamSq7uv8XOZmgeiSk3qsQPGQ
x2d4nP615yb2LiPXuBOhBCtKztA9owhnJjOMbLhhlbiYIsf5ON88CX7OTWSOztNzXAonaYMYwWM1
ZA2KbJQqm4WWsC4czTmSPAk8O7Aq7jXl+/kc4ztkE6KIw2t1uZpEAdMAo0JENKWPZsSjCRpaMCVp
cdN4khusHnFz2t8yIjMe1ARFn3xwEn5DTEzp0GX4KXZBIkoIfMi123OyA8ge559SWrQV5ufjnpEt
EefMdhr+HM2wjZmiyAn+IOjav/UO6xWeEcaFaluTR9po2LDOg5X/JOSHOY9UDzKiO5fh0TgGYjV1
lwXuN8wVFELFmpQpYKOxCd67mDJDtRDKLM9u0KONvRBreroDv/YsZm5h3RGpXheqQECb7n/Kh5IS
p2EPr3Qcx6AKGSVCHVYABZYvNpKE2V2Y2KJt7L1s1PEoKsYFkzo/YCNqa0pxKsVxBu4W3JL3eUkA
TZ3M/mcpEqnL3+CWlFK0l6XWSmTPRLwCxHHmMKwD+3lSANqFYACMNE9+iRVo9lHvXTbTA64/Dr08
u7fJuH14kzVRaAOnCYw2SL+JnJJUlSj57Em3UDlD4YLwo/SDWzayjh4iMl3YmcADOAuafwDeK6i0
ZA6BJOxvOJ6y6opTksGJlQAPePOjF83ikg0nxjfAIGqRJo0cwVNHcMYrp05zZmzo6R1sa+Bm7Fco
fCEH921nRrEAEPmEfrQFQbiG2/9yVz1uMMUZgW79e+QBlMvVn4zemWipeM3hIYYzJ32GNwb6i2bD
6Wcrm1LlBie9epDyto5VuEnHwKH3kJdD4oHHz2iEZtpS1hV3JGTtk+hcCKjDuKCR+Xnn7VX1jn3S
uVpPys9QHvMN9Sj87Kni6VcHiOsGQuKg6Qiw1Ratrv/l9ppilICdR0CZDps85tMWWcgCat4Cf4yE
taGAFLDNkFlhU+7H0iDDrtDZhSUROPYyyU+kCsNqP1F1KKeA8qefyhI9oolxRe/CA4NiTNlKpRt5
F7LZ/pDdfJrGncGf9gv/mdDtek+hBB5hvTseS5JB3TvEuUpNV4naPN9Yzgpr/tiLZkv19nLJXVUZ
KNFcm6f2nxm7xr6yn+V5DyIXoXB7N4dpdJDaIiMQvXWarx5UdvOwCkeom/zcmzfhbz5XAd952xOh
eIuGZ1c3pNHOuTSVVDrs7xRkhEL9rEBvS8lJJqI0KQK0N69hntSUrDgaT0kh/mt6yAeAURf6+hlg
j7pEJnmsCKaG4q4SDD3qK0y2tVht2r7IxXA+/0kF9B79Ck25KNGj2UWo4AveizW7Z7lu7lHeqwRM
KYWHxcBhvanAIpzv91vS+qyihNfO+N89EDoO+Gdr+VeP2WSPkYtYk8CwswPlxruRpBTTTkUNxj7Q
bf6pnIdJFbmzFKjsgqrsCjhV28JNYEvIM0PjxGw2G3C62+WF+zf9EyNLhQ9FtqwqQc97c0oKN3W4
cZo9gNZOuSlBKzhAHWyiP4e+yLaQkcLdnHZb4DN87++ELneNK55NhIEBlBm1po+hnwzTNi9wkxNn
RewRuEEyMZjmZppNeCX2Y8Aawil4+uK5GtwfLm593YM3iwoeeyD6bESY1IRsq8IB0Rawto3msKHM
2OsWQb9f8t6jfnDkJPKirDM2r3EvSQaDAvecMNGnBmm+BLLixDdSzy36hEtsOkIgtz9h5FjO3TQ0
lJAkuzbG5S3Yqo8/houSCnYH12llt00puFWc8fEszWcco3UY4gXpC0Qvccr00TT0qhPPMLGG06Gz
uYjENY/qei2ri+1PN+vSgb7KutJB69oeFXQi3XkipcqKp+PCluGG086GurkafsNuu3h88I3OHGf0
7M+nzBTMJUTO126fNKYKKyZmQdU57ucvljSIDcBTtj7Vti+WEqX6ViLMaaL4XjM+xdkWiYsn00BP
5lfqEES19SGYQ8IivF32kOgJ77KS+j4sA62yxyFyXPPmlTEzOCeJv5F2F3b4LxzUS54oWk0HBfQ0
qJnLtUIX8Hn51CbwP2z5ieha0jUUwOj8z+yE1dZNmGiRNt4L71TjDmWXpxMiGTMmzSSkNRNSKmbS
YxnYP2+7gLS/Z9tfO5tTVjNfrJ03B1969u4OmaCORkQaPruN499K6Ly7187+4ZzrvB+8LnMa55Ba
sdwRDl5z8oUCIfr3l4habnRFSNMmmPuurRtV/NwsWK42ZgAADFmxfbgaHmaWmTAFGktZqjFmoXIm
sjz2ekW4WLMvkiCsDOIRF8uc6UzYsf0o9QGOVb1LLogQ2wb31mozdPXP9hwyqkAbxW6JrydOmmfq
+tQ2aRWR4gUIDQnQ0rC1IYu/gIlHOl1rIaPovNFd5TiR/B8mLxm1IiRIKOkZOLly8tTLc2lI6ghe
jfCsxMiUP+U+qH4rUqiQjTYn809ywq5jZWZsZeL5kFaK/7VTnvm+KiaYz6DzFVsVDDM9aCSwqJXk
kRW30X4nBUP1R4m4idAiEyVNKqlD3owBivOLi0i8D25/S3Lru1YUBRzL/D7zhFRV8ruk0/cCfbYc
iXiLsAnNPxipSX+A88hjH7rug4Mqw8zGNmdhxDyALLQL56bHaNU37Jfa17nco36vjxkfnhOcUCbM
yX3dkrMbu++ZYuo185vOkpOO/3EOG59ELTqxmwajzXCzjj4KyqLlEoUqD23RUVKwVuHbP17UruDR
D5atFoQXy2f8yXL/8JrYHNCJcm7vZeE5D9q6wxsBIooAXEB/oirG3scbqWSQlAAT728+i5Rp4ZXU
Dis3cyNF8wSeSkOhb9B1ROYwUW/RW56Exp7MxdUqEknhLzfiIX/m69Y5SnZb+b+ZfaYKffshEHwy
bHIf7Qg8tBboeVQPXewc0pFTpkBaYxSTCwzUarnyqbvURyHsRVpHzwmUqnqbj4MXKuiwT514sOEe
4EnNO9lU+sGVQ5Ut/k5R2hgYi5GwqEj2orC5SKUUL2hdZR+3z342vyZ+NOF1rhRVg4VNmLQ/uABg
lDRUtxsWxxQ9exwHfWxLuJpzOjKcHNOjcGf8Ld3PDPgQ9bT1envuXo/mAxCGKWG1CWq/Jkbkuabv
CgKGao/YPIvrQd1eaBPFipL271DeygjZ98GKEetn9f/GIynO7+yzF2OfwRuyBCeb45qB3znD8Mk5
DHXgDgQdy3mUJypaGSeD+etVlOGMBSLDA10jyulgpnU5rWTF5NBCElfBkAX1x+V27gr/QyAkhz8u
Fnaw2MRx5mYUZ6nVmFf37+rI3Tlpa7xcAWjIQxm5bZTkiKVi0F4Tr6ABN1RjxW6JmqoMwFwcUj+u
EPphSA8YQvP07KcVcQ/F1uAJZM+3Xst139w9jN3Gkt7Q4yr8yG4oIheZiSIjkHM9FXKgCHsSCngc
BDlro+hgeWjNI0hyr0vSB8yFj4mfBaVnAJhkUcdv0BYYvzGhShmUJSp9LQotggf4VpzsZWs57IC5
fn9u4IlxDsulMY03qd8kpaEfnMporzkfyGRBhTH8HUTEPFXbTdSOsqTx0v0pGKTGuy7nsmGLwfAD
yTkO6iWeqDQu7O56OC6As1WnbMx0uieAyggNo4+f745cxzIoWE+Y49azN8mi3N+INeWbvx5BUNSL
V7wCX7zSLpImsOOakp31Hn/pw5R+ztYrCFceCbIpKeWeLFdjoA1MMXEmN1h6nGhys9GShSPub+I9
rMAqiiEaozS4fNKShhOaoOAnQlfvYp370QoABGGoV/felWSuzUg/p9AohYURbQU8d9tBVWt9huZo
YelTgJeYeDSTjWhp5jK6W/RFYtSUeXeThCAsIFXS9bHSqJXOYDuo0aXnBubngp+zEj8rVVLgBzrn
BptBLb256LwWd9gED/bt8ZBED1NIZ/pvZgGlP5Ej6RYR05GMRJG2UKdmipMk3tlBjLdzupaPS4b8
Qxhf2Z2Obf/33E1TjnNSId4DHGt/Fl3O1WPvcZMy6vpW23+3Gk6ip0f0Pn0AOxHXI1nTr0I783+9
/RNTnhR4n5hsX1sJ7Sk/31ssglxEPWA5dliOAbAZ3o740xq3/aVKG9MOdUVK/i7uHyX4IAiQO7/x
M/IArFctmBXr7sOvIdGh2WXPLARfvNb18wnHDaK5gZPaS8DaqVbnb4v9FgbYPaGSauOntDmHMxt7
sBuEbX0Kzfiu0Wdi2oXLCSskmw7AgwffnkXVZ3r4p1wrpPQC0tg7kmm4Gvk0C7WNhefDQZI7EVbO
Biwsp5J0EF+nXA8HIemUO95+Oxvc4OR1Igl3Cq0HMzKH/M68ba3aDx2QOn4BofrxpUO0t/6jE6rj
j1FbfCx+heVDc3R7g/qdE2bxNeKvBpRre8Z+Kv17eg7GnB2vKwx/bxH3yRfrAQFYSBs9bjjdd7hu
9Yieknsi5RcICI1Rq08VV/LroRlVgZDd8kjxNMDQ/Uk7NPArkUIexRPLIRr2zcjQjcuq1r+zVukw
mpgLS3nuQTnQ3p4nokcgHol0j0thbkJU39Tq7xUVFj9r0RNq0pybZ26o/ra99+r2okEmswONRbcb
kcYZ/Gf9rAsRZxCC7Sk0inpKpUwrqGRTmQmzSHRuB2bue6FTbyeTeFEXY3WHeZ2v4uuhfUudeFkf
CnJqLPaD/HdYXJLFE8In+RbuinxAu0yFcP0OSiaDStRlVF9oh7JLMgbRgEtjUPM2pfBI905Vb/h+
SqrB63iQVZYsuT19vmn8pzZ7BPg/qEHGDUIklXg88T7ab/4F2pkbCBJ/U1pu+nj5wsXFp0j54GMS
je4qmXs+dvE64cJa5/VVyRKxtyOXZHldSPVlLQyQJDHIUzhmwCF48WvcZxA6XD1Cy2v252a55DJO
OrSWJfTsro6T/wSq9vFtlcUL/UZW5JDyqo+CqFqD14gUNjGpYdXWaaQwuydCGjYv9sghi3X/fvZP
Ih7Y0Derj6QLyMr0tFrNlq2WEVxoLHvC+5Sml3dnYUQlFjXKtdWOpodiji41D4MrGA2Pul5KZtb3
LwJmBy3K1it8Y93koAjVKb4ELQ5ccFliztebDPmw49F3iW8JdbWQBlp7/LIz9wEAemExS51ghi49
LONJN6va1aOgmt1Lkxmlu2PCbziuL2SJ0dgbigk7pVbQt8xj4WA+JSbhxj+Uw4MVSgpzjCE0SBCe
w+8dRjrPyYY5aNuJ9KpsQ7PF3xlXXl77zCde+DBQ4t06X97Yf6K1uFaTivCZfNM0+Rq6NoXzZM4h
Gz5dl8oxdd/aNbj3WuHd6yk7mQHo4mtpR6gA0AC/0PpxOKGBWRdy6Hdg5oUm0Ts9nPz9UqbzILLw
1DZWdVqLlWLCZBmsmAcf2NHbyjU5cuvWm3+EsIaV8MvvijJUou3nxHKsCIozORZ/v+A+R5ZnBJrZ
isWU0JX8LeamcarAjUjYn+2+PNJlyGboS2XmVHphkgfwY3HiSHBsxQQeyVtTvt4PoUBSrK4XlbaT
EJbJ30+6WuWM4zkCTxhxyoKjeam9SHKvutHAL1U9NCSqmkNl0EdNiQPjK4QPgbAkDXO9RezKZUtn
9FNfR67XxxcqiiRPsz0u535h4MGWvpR0V/N2t8SyE4j4frtjicSK016OONbjQsgGKNPp0oHYcIyf
kGJ24Gy3ERmliOGQ64RSoIFRwbTq4mJ2gGwgNUVgybkUjoP1/Ba+MFKvpQoaVAAP21clVYafDs1o
Z41KWsIPlFNYeqZVIywa/mnR2zHKk4SLYVwOKUHOWvjurWfY2yCKGjnKAkV08hxPXF5FX9+xqD2K
A8SFKGANnm35aFiuHNUtRfAVVT2CH0EC5QC4sNLT3cexUgNo734t9LXuK/iDRSIDLVZtXw96zl0V
OJ6KLRuoVTtlhydQpB6G5oKxwCmDz+Q++LPDIrGooLzawMNExoRuYUIVuZUXaFvlBW+CVvqDMErP
NDVexDpC4aUkIbmJ9AOuac0CPcVk5Wvt4dzN/E57APVZ2ZEibumPpC2B1FcwIIE4s9Yro/2A5vqC
KBxRNAR08qhBinGrDhjchDIyDPlsrnNVkGSAiBIsgczz2LqWWrizT8VUc82Mb+dDxlabKsRYOJ1I
h18zRmHR1Wp7AbWSorGNnIyT1c/YET92NqcpVCKOlREJ5lgpBJbcn7U15nuChKvxkMUuxbC4t2y7
HE6KQUFEENs1/BjLOqIPOeeMMiWkxEqKYkInYdx0tLWk8q1vgx21Eauc7zhdN1fxGw7y/srkA83L
6o82B91CuKdRP+ufvuCYNoyVCnpOjf/F2nfH5a673fW5352v0MvM4H6oE5PHQ/Nr6kqYorss+d47
XnqWumgiPZqN4i1TchchWWgnVccnynQ1nBxWxyeq+vsHKKh9Uwsaoav7cTDBE3aSI+gyp0kkvVKf
Ky+o9xKaG+cKDo4HzSKfNh34nb1HWbgMFWqtydIzG3Uzrl6Yqv6Gfc4On8JCrNNSqDaceddquJAo
76HTQWdRY4vsMp0rR+bSi6vXkf+WfjVlu2958Jp17AlTEwgs70t9iBLLBNetnYHEwVDT7lZSa3D3
RkmafXVrj2O3rMp7GHsfqHWl2fpN5TgdiXC4NnUhjgnU1fB4beNgjADdhvXilVjpI61HuinQXKHL
DiXtvwuydsjaRo3ErubXaQDah1XzsFfTKZIVg+AOeXnH6GfDMZ/UskjSRGX6yjolc8xzfNTfnvUo
P1hpuNyTIqPJ/ew6lnLqvJ9e6GUAttDB0yP+C/WHVth4Tv6Mct6Dmku4Txfsf2/0bJ1QBBlGrcOb
4Ply0m4H+YffJARz5gxRmAz9jEcKDqssw4h3EuMKPMhzWG4zRTciY+7F/U+9UKvh/xXuayOpaewO
3qbwVOh7f0Ox5lTiQXOjnqk+V1shSrRpQIj1OUK2N7YYZcjG+jBIKeBiFzoF9Z5+6PAovk4WUSkj
m+Z7i05HT9MZbOjnkggNdXoebd0camKxRIXbFqVIfdgbBvPE61p9lc2Mhbw8RDGjteoApf/8orIX
Q9juCR8WcWsEwTH8G6+w+KeWad6BeHECht9ddGS6CIkVnMVt+vwj4PI0THMDJsD8gpdju6BHdeyi
MXM8z0JwE0DwewNX0YFuiC3sG4JMTYhHzi2p5ZmPXLLqdOJ93VqjU+2To5hi3+ANZLx49YYkriK9
Fd7JKx3yxs7Qw9Um+Yr5krIQVbvdYis/D7GMvm+Ky+d7V8UODAHvYWVgYCDgH/CzSkIT5u//Dz9x
g2djxMSjsgGigIGMcKnNQCxZZM7lsAM3X7JV9DdBVId7SH76fNTyU7f4KGz/bltswdtCSr8IlleA
7QGbOq8pmcAy9AK7FBSE6xDoGl0TpBsxUDgcoYwwPOBnu+yJ46vGl5oM7DYQZ08DAicu5pn0fbF9
w5co/jarV8+aqd/sH0t2jCk0lSX3O0rnOUrrtXbMdnYps0r3a8t5KV1RCW72pg+sxOkCIKTNZjR7
QDToj8XLZALSaWz9Ug6a14GEwDx8JuXH9rnRubG2ljabETt6H2bhpTYpfNhj4vRfps3s1yeU3Q9m
db0oQJAZI10YZPGa5Hr9DuSYNX8N427COfWxCNH4EQgJRbhcm6HqbOqd9wim9XfAEcj1Tlgf1WIK
omv5KOtdgm0Pa7fHY+tzptbfw7+1v5s1+0wyfWOSqa2389k4vDGWxX3yR+Wf5h/D0c2nqSFkS3LO
v+jd20MugjCeS4ofb2sex5oaVqqMSK6mEGHDfnjIFYxvOkYarvmuSCjY+oUSp7OFTFxkP454UJ+6
opDe06eOf7aShZLzgjYoRoOocTxDaCrBuLUl11E7PdCPfrdDNspx/R0B3deQP78rHchQlv3VgZm1
8cUXgmVfod5FD4fufdIYOweDXOeiYuMn9ouiUUPBHDskONI3qBS7pZGlYFJ8XisUFPm0kbqCgTFJ
3jOSJk7WBgTabgj8opOl80R8lfcQVNCPvBZMzn3gdFwIly7BFpmpuA3tB1jZD/oGASXPfvzfVBkv
1feiZQSkgBWGRouVCUNtipMCbcpRpJLUr7XqCLwzOZnHrbPlPWMVEwXN49OfKX7PFI5VjABWZB7k
A3q+f7In1YrYK+GGc2iDH74AUPko3d/rqTRdmL6yTLYfOkT0dC2YZgIfgZ2ojNBVAWTN1g4Yd2yo
/wCEg7DrI9AleVoJ2ZpDrKcItCG837SZBpunuhysNCXqj+apaYq/qlhR555pDBcaAHC0LMixAILV
UMRmQ6TJdsALsUG9ectnkWTTgsm0sJd0eNRlL999u+7EzA4UCwAtw18SU8FLqGOYZraVYZjC7O+a
pQi/2Kg8XR8PGTu0xUS8kHSmuY4d/0YVfi23HVyo1jlkKhHTH0KO/iqvqLRABirtq/Qu4/xjZTyj
+hynH89fZWLf/lpnlvYpaNyvLK/pD1dJoy7ya9Gbr6LGe0sTCEJPJMMvlQiTFlef7e9wmiRf7VEu
v/9efVCijno2ox3OF6LZyn6ftErXN1gg7Sqnuz2kR4nUFELSQk/0eYeq3Pys+rGQIZuEB+nWIw4x
Zs9l6zTWxO8dll+cKRF8/lC4K6EoJkjRtbCSjKXu5vJKQOhtG45gZjAJx6jOSEsJb3st6aBiqoJl
nO6WqAMV8X4YzFauBnUf29y8ozwkt8e+AmQaQrSZaVwMY2/268KFK5d7mCoFaZYb83GZ+mSHdb/v
nKcO+5xpyJSQatz2awxWXjh77xsF7W1rscTmHzfKiT9JQlg4a+T5FbJ4lIEFZZS1nfW8tIX1M4iW
dzsdmQ83UBMQ7UjlcGvQgFIAiQLkTBBryi/ogT3l45/kqs7wW+STXrOgYsjFbtgeyHB99+NrqqRl
IWaSQbY97nG7isOzAEO94Dtb6EAaSxJmIyxN9bfGlSUtBy8+ZMTeVPoHjTis+WafmWHEjNHpAzf+
sYK+dqIBvTTcgirv4xJGXJCcpL461qLDAmQWnoxfaERXcbMVhs2gRZMeZEV7ivxi0tEtL+EXnpbT
JrBHlLu4lUfa57okgeRtRuKSWFo11MpBBjMFc0nL+IRwlpfsW1NZ2p2Zg2LBt6Sg78Kc28Wrm31t
q4AUoSWk2/ggYwAz3F0yFJzfDipQT0W0vDx2dVCmjQTF+bo8msZEdLBKKEo3OdDfkVyipM8MpiIK
Q2sbXAejbvmFVk/1fIZ4VplOO5t6QGy1uZxm2Px6EzkfoS15Mi1PZEtAz0Rhe4Mn0NjMW1IpimNT
jD2l7NYissiMVeM0EOh7YNLEwKxIf9I8/zdEgyjFZwQKfCGPAgCxIjYHuVAg/xOLORzB+BAmjOAH
1/Xdu3Bxsw//IXk7JQKjfMvErv9Jd7pff7R1pltIG8SwuAsZaJw6/9PjI2WAxrieafJwI5xIDzpV
xmMepvs8jQivPBUlaucQ/rh2DoA7Apo0Wii/iA+9Xta1phB7MjjGdODW8lWaD7nVGdM776CkvELZ
531RmxyOIW1c9nPKb1YaDflOjsaLI3IzVVb2GPqL7RSNgfeKzEIuo9PRHLOqUsj5U1XTN7xSzket
u4AmEXltVN84xNn/ErnaT0yRXgpwXndxL1b3YfVQqa+0ZH8EFEH3DHw4Cqjc8Zi3KA+F7fXZlbv/
rIsV/8/MS0SzOfi+OQiBWvvRxL6ocI4YKjVxycyFVzuxC1S1cdgFSow8EPz44iAo4jWiug5yo3aR
KrUbJC1SuC5vP16Yr6yqLaJW7Ymushn1LHwa/TFGlE83SzFGvXdCav7C1EwledJri4M/v6QPpJIL
5KmP8Q5T8D+7H68pJgy5+qVYPlTrNpPAjf0a4bGFVxgXulVvNG0ubhTvvGI/+9UpmD1B2uThjicI
V80OPYo6SU4kMzQJzRDD75MuWeH5tRmXEJW6nTahlSHV2OpQEHmh50WTYslxbRK/TF9q8piHtKgc
M+xCOTu18fkvUJW2kHK9FQZwnzfOT+2f1W8lbFX8ENxAXbiTKlcKKblfC7c9rgtpyiSg2SnBCLu5
O1PascGy1Z1qxF1Gmvy9s8Igk7ERV8N47FA8FpXoj5+e2PEdaAbB6O1yRjZLJ3Y1S5VTq4PAJoY5
u8qJKwZKrvR3kJ7f+bYtitL4lEdKFx7vwKo3zwx9zKK7VR2LuDkMUD0/NDcdi5/pXmfwhiWA3G4G
q52vMkikyyagj+7ufsbRE2ZCUUqK9tceQO/u44fSq7ugSHmk48yV98ED3PGE5jkyTRJblyjwTLE+
8GajtIJkKoP33LVtreLJ8fgND0FF7C670rI1WC3SBx0Oadm03xShXhbYE7W5K7KuAiDmTgnAwSsG
QM81LvoKzTCGaAd8zabMwSD1d69ymJBO++I/mmBmDJ7lDvUZzM+mbm22t0nHk2nlmc3w4CvTf7Jp
b/UN31rvWVYYctlyAe/vPieq8pvVXDjE96E431Sq4z8x9RY/9RTcwqxMtkwXpBz4IQ76/0gSaUC/
tl1lYKmN73jHTFNmYbkPigIQm06ze6qtV1Fc4rVj9JRb03p3wxEvWcaVUjC+Rftv4Vjy2QxQDxgU
ixnaOdVxld6aS5ftyxBg+XAiefhaUuMb3+GRxVJDxdv37eIzfBK8/T3I3Lh7XBUfYJgLa2CLEYz/
6oPckp/i6eo73a/plfgq9z9xr36vPDpqMZXs2MC1bOAcTdySK+t07696PTcBodDTfq5Qsjn6RDpC
4USnyztw84yKWsHBgUpBU6NY+a2W1F3Hv6bbean0lAGRziyP2LudoXZ1MKKDsjnKSyqPZ0zhgoNL
EZaVxRtAKDPNZFmfNcpCxmTXxIB2lCNl3r3p9zWP80zw6TUvGFB48LApI/rww7o/MMbNEU638vDr
MMWEVvL8kOOa97jiW1F6xzhU69JrSsTy0jxlJX9wqnSzTHRzcBFzkiJfb63zETg9uUI2xsLbtB1h
oa4GmvZY5xynpLihB+HkHYyVBwIRZC6dEFntsh6KvJmdPeDeeurc8RqMvfQKNVkVuVOEgv0wZ8jD
HRboL/f3qfKi7RUM8tVcTAGi2IuMcgP4McbC0GlRYGw2EIf7uiArcvTygPa0YgyfUZG35wHsUtrV
WW1jal5IKlg6f0vkSbm351m381HyfJQOntIH3CwjHxNX4LhmrGEree9k4f0BHz2/f17n8rDo39lb
jHAxF1cJ1srfxzAWknqwxf6Jk7p2C2xyoneyw93QUsPebSurWrRT1+UkuSm4kWCWim80NHUYs09I
Aflj69BQ3TAEIXd0QRXsTKeYs5wiDCsPNqAEMNzqdWWKVC7vj5KsVxT5bHKgtX2kgw+VAYpHHxJn
PGZ1Y7aDDY99BDq88ENDPWH66ltqHZ2q+yLGNNDZGbmIreh5L/Hj2xP8Ig1c10dwVyTSDNaiMVo6
35o8SShhykdOfFMvuNHoixGkImV1hNZpiErQNJHJW+H4IWUCao6AKqsYafVamS4mSzY63E7xMqRD
EKNHnUzvZmlbLFbU62lPJ/egAikPoi9QfW0muasRON6Ed53JHIE6wXjivOOvQMgmfVVTyuKTH0YN
C/VSfqI0ZeBKqJz8O1wu2jHMeokMq10O7dr26fOnv5NNgprAEbpnVpMmIDsgzEobveRWIqO4nBQQ
1t/fDt0McarblwW0HGbXFLFf5ceNLKwXmTY1seGeC7SskOVkq+X06mlPCq6m67sHwJcccBLkDCi0
qM3I0tprkPCoRJ/rglPgpyt3zCZceBj+evzOxC04yl/Df+luir3jqbYUx65A8wVQOVYpMXJi3F+1
ERjetGmSsFFGmJ6K/hBFJkwMbO5cntH2unLK5/yU9/EWyvDqVMuZRGmH9CICV86Q3A4g6nXLK5IM
xjN3C6PX36ASUna5LH1XgQ5cUQ6VTetc9EILD59VVqCk8n/VeNe1gotlHXbRdU8mL47BqmJ70EgF
1//prnj64egxpqLUSwZws3tQPoPKjoxPL74X7MZ0A/06gmqss8Zs2+q0u9vY1a5NwTtDdkFdB5tE
5pTJvM0+KvPlMtnVxOnj1J88F9Q/1QV/iIWQhFJHguGDYmoR/ld4QJ1/CcKAi4HcqO+JvHjqOKjo
BfMngV8jaDq2YTpa7tqka439smgytkJltpljwoIsnv1e20XVV7kzfHu5wqiOZUfjukfnvoXZ5CQg
N5s7SbexbaCO3leh4wwIFZWppWhZpyfRUP0D2B0AztZajReMxKg9z8mISP8zmlpVpPLQPyMBRIC9
kKnhBwPW4irNgb7iqAfHd633QiU4F9FC9zt0bZMjycq3mgqwYlXNKvTq8OHx43RTeveZOdioUldC
s+daNd4AYXkhCtgRGNNXceW2sPLUzziV6VKce5iI+b/jkCqZE2so2w/D26h3VeY3+fuSEBGZhcth
d8qSnNWv/S7mMHDqNEFU9AT+1mOJTtkjS7h9y3oYnBkySmLBmyKeOfi3zerXRA8X/RdaTkJXV/5S
A1tpei0/4gKDmh1z2NDN19nIQt2tTU4w7FYEdx7fMD4quQI4sKG8v+ID4QUUr14FNwGoJ9SIcjod
DJgQbXSwghS4RlA1bNvCt9AhfQ6yn7O19saMzzidkhtYrcGUYGseovp93L38i9NEa4qzmYYqcAJJ
XLBWJG4NhJYokJK/KBI4gXFn6Hl0zqCPA5hgxQLPuKF1oq6ih4Ul4YK8f9SgOFlKI/yNhQmKpqt6
gwYKeVB7743twnfPmbMpX7PHZKdg5SkAcFpz08wpQLxezV+m+67QuW+9X5G7jlwkKzJ4gOudqyjA
cFeoSJ9EQHXIoeX4zBn8A0BoYAtD5Nk1ZTZJU3PFwhe1saK6+YtADq4Ynb/cCNsNj+HsFTLWKJOd
UwirzuLMcWHWVaHxsGGnr+MN8aGot67ACRECbFiUc/poRsTIk2PIrxhv2izOAouEd1hRanaTWZOq
tTactZZ1h7uQseiETk0iGXkBc7jv3phmtq1E9En1hze+ZYnC/OSen6iIauwuolyDk84a7IF9IhpB
1UFYs8UES3fksTVS+eebYPdhedoY+4xSdaknj+dg9tOZGzsXE5E9BrgC8KSPMfCnkrDYA2su7APl
WfEvutJFYO3KbmIaoJxLIS8UMkW//OdzDIx5Tmbk/4s8iAUhJ7DqLby4Kulo1h8tBCZie25q8O75
ITweoHZrBcbZiPTiL+kENRyAGauMeu1HrUs30a8eUlUBG9ry+g2r8b8lFjHnn4L3P7L40apmokCl
4AMhPtUBe8xcqVyq8KgOE5TVc0XBVwxG/RMvGvuvpsuY/Tn3LvumnHN8P1FEIf0WZzr2+96Zm9F9
ugpNNN3gf+buu2JSRntKx3q09omeUP7Ybo7kRYy03ViiurzdC770HBShYzNvHNUkQ3QzFtdI07pq
PPywVDzMtTwoU2fhN1s0LNjS/GufVi1qJQA4WGsC4BdhOBdGQU8FxNu9mmc90D4Nt+iJbLNN1le9
fThswdI883vVOEml5TDjYYDLQI4BqZzYgsgCXKmHT+Ut5Dmw+nXB3PzaQTMoFaZb6ZgDd/k7y3vS
8gud4GcdlLkXMRxM8PHrkkGF2OcpVWsvXXl3rKRXALvvE5h84S3E3STselNly57BfScgoGotnk/I
NKwMS5SDSrmHl2eAdjlb//KxHffLTOVdILsze9lwDGCWobkAQ5nm2L2YuOQn7cADC76cK4iDMget
ClWjFYx2nj4P7yDUsLQRXkzMaz+i9rjfXp+i6ljDdi+DnAchc1r/noqqw1iu75rbvUQXlv29ln7O
AwHXZIZ08fGJEXSON7ZFoyDxFD3dK0Zabi5wulTTQ/IDuP/FqEnAfFxtW+BPw/Dh4FSStuUQTukg
CyJvw92C1uhHFay59/MCQq8S46Vk4R5/Kra7evMZYtprt+aQNUSxp//QST6q/oPS8PV85sDSc2Tt
OkU27Gg4QjNkbvUK3r5eiG5PI1Lcsun18uhjp++tt5mp1Eh28fKVi1T44/QAXZoupxA6CpW0vCAw
HKPWfnDaYeKzPE2b8si4RlbYkEYC8hWtoMv3bjULU+DFaB0OO24nZxm4QepvRJOWidWC/iu08X+F
wq6rcoOVaOa+rGaCSDht8gKcGcCuZq1MThCBGOy3yJ4aYsTysA9djrZTnpZW2gDeXvn/xtnQAcPW
r4sHDsOu/Cf/ByjwSop0CoGw1Tq/wl/v45eYvqbrDftJ6K065bCiFXDehBO4u9rWSbTemURe/FHZ
wgR+DC+xb8X6RjdFlQpgtEoD4EaWNsXDjxYpze8AjhvGpj175RrDU8TUyUm/cnvkVB8kZb7+ai8t
zNi5p9JUFEo/ax9H3Gx9qjimOsc0PpsGugccZSGvjL7tnCNjSO9xTFMD9iyLcNzWYdiZxK8lrDPO
j6YwzVUEdxY66vlBNVSaQeNmBfJjynT43V9NXVTI3hjk35qNOh5000VVD0nWn8wc4WSAfQt8MhxY
brRIzmckQe6ZKHGQ+leRbimmpp+y4MYc5v9JePtEO4FjzIggAbTrof4oktkrjIGDEw7kvDxd5yyL
EBmvHl4JHkjT06UWukTEiJVkiIf4wY3L1EtrxZ7v0DRAkQI3B+TUiD2mGTaGE2x2dNMrHlU51Ii0
Ja8Qr9Fg5IFEtIXo9D8Lc95k11aL3LMnfKSnEos4kwJxlNyFLw/0n9jp0Aq+xqUV6c7Dbek4NmfL
0DRCiLbUYSQU4fUtvMtbVGiIO15LFuiGmX+sIDRsf/VcNgvoZ196id3HmvQdBEriA+oW6F6cPESG
io2pQRU90J/7EvOs7HfRmJTNBoAYJ6vKa6CJFVJQhM3kyRzZeJfbQBGjpbwyEm19/0Rwiv1p6qCd
gVrHop6QJ9Ji9YxTwCqbYkCFqVZJ3tyze4xyzAALgcF4O8e3OeBe+9dGzW00v9VoMJhjzgvTjz2k
jfKuUYLdDiOCuin8Ftb4HCqRDqjGF5wOvldJQYMOKVDziaKDuhtIwXmCXmsjbujIMwry/1l5Pup/
sRVm655JdkfcUoHGAT23namSs+4O7pXn0wLDBNIEriyU44UinK5h5uQtA50n1ZPhJqdBcJ2eB0pX
dpIJNGd/KlzNUyTIkyuL0Ktcx64uo6Xyej9VvpwjbLJLfh59GSoEYW3uleJ5GhqYBjsrXgWJQGRg
xJCu9vIJeu06UojzMx9xuDaVuQZDWdC3bA+/QUA0D1eMzNe23xuEn5pmF9NFZE32nrXdKrlQen26
jDcgSoGoqIzrTZe5gGNKEOeW1UxMep/hbna5IhXDEHrWFtokASUVi5JIQraz9Dy2jvjhXMFEdkIG
A/gLEFkTCvYVrJ4W+F9IdVLa35dKChmGA2cmeaSiZx5URv0CG3JdJPl+JlRd+t/mb/PC8gjuTsnw
3fSJHAraLZDcCz+ByTNmQ0RGVEvrmT0OlYesTH3qZwjzBt8QOWp/Zr+24mphi1cZyoxSbzMvCqcR
oNyn9eQOJJ55Y8qjiKrRq/UayJa0ZD1VVu56j3YDrihA9AcvqwLeOOIWYIEgFCDne00E2HtO5LIg
STwCqdReLUWOSMNnK9AwGxSHLM5DetZi9Zk4P0QQ6UjCffslKYkOrn8TwcltCXmZpMq+HKJTH8jF
Zc0GJqDpe1EKFmxub8SMs5uw+Ep7kykIyR22v5U3ppemP6U8C48kALmfIxSbDyWP/lPg+CAqVDF2
jQmVBHTPz+2KhQTbmB+FJil+K7je1DMf3bEN0d5WZWyDlp+bpDOZFNeqf5af94xgARYK8U76lZQq
0LO5fQw4+RacAut+on85/WDY6MOY3m1hCYZiHYlYtHeNPSQTu+fqNqz9TO/5UcsE+lS5k8ZjahB7
8jg47szmlLILl+6YY2Pq8en2lExSeiyFN4yNitQyP8Bi7EA8GHLWDaR1z5MU7dPantErzGkqA5s4
r+Q0qwqPftrwyCn3ZhfRLBCZ0Kq1i3yNQbUV52xJZoTRUywSZsT/eS8PEmjhZj7j4okoVWMiZ4Nd
r+LaeH2yj87jxoRLTIBSlLU5dVWL6SoQwGQlUkfZssLvQMIuKbTp2lZh1wYXcQ7rUZrasY1JuW2e
uLLoKk2Oz9Jim66h3RXWkpIXjNdjTbmXQc+pOg1UEwljS3x1WnW8aKDRBaUww3Gc9Fy7s7F4yRxY
bM6Oo7HhwD852BtzvkryN0mgz+th5w2q4CDjmzhEXI8U+N/QnytDbqArxyovN9aH2y2o5HC5f4Sp
RkYIKqbgMrVht/MIZegf/dz6p1VZpDtsyDynhe54ccV59HIDeO91gvnIb5EoBTWf6f5ZKKMltom2
wvVs1RSImGAEgAyk47hR9kymHzPV5+j94L3lF/RPbunx5qlEt1XGa6AY+ujMXUeG3zCJ2VUVQDO9
1wKIXQaTXL4H2bx0J1wvMa9mHDa/VEHNMYHPd9PhZmlkL8y6heIjWh2FDuRKwZsVCvQ2gBwaIhfO
/F7ZRBdJjJZ5KO4L7roD3VTC/wleNDG2qrrVnpXq0B2RcubEpEV3Qp9gkDNxR7ziPM5nv+HoZ6Lv
AGmS7L4njSFTCAbbfSSuh9v/sZl3RZqXRnS0c/x4XdkzcQaJo+plqIdCYnvGA//ypyneUW46WeYL
P1cA8xP5MvBPA8bpfFH9gTpaQzXS84Ac0R9TjNlipZjVmKr5iWz0NXRHcCndH62nAaeJRmhoi3ma
/d+WjNAttp5uOC/+hpHLjCe73iHrIcC8PY15zVkgb0hWM4GHxF4vW/SiFHDjN71aV1KD0OrCqpFs
ecU+kUSe2NPR2qLAhi5Ch8GgPMgVDP0bAkQTCEY33nQLwdYeeKtjE2yldss4/06Lzhi8mTzNNLoP
qBnliORYhUBTTvYojju4NNL1ePqf4ytQ/brM8SyQzdTcgBJA/6DFf48KBtShzky9PXFAyQ9ACg3e
58o4Efq32svpTDSqI9m9iNwSXryiRA9RxNp2Onyg6376jB8JVB/QLhYvCLNKHFrbomofmWhn95un
al56OIT1AJ4AT3mQVoeh3tQ6XYQIh34rNlG6g9IMbOL5WPefOPTDHnrX8a0amRncipt4lFSeCC2N
4I6TBA6LralYikrdJ4WidKa/vp4KKSOKORgSba/qkGfNwkz3B7xpdzlPMqSmbCjf/XjX6N0Z5Hf5
uzDkJmczR3yhOBuaBEdaJTnS5xjaBbja/fUuq96oMWFB/GcDXNfPuumYfqfiw1kL0NX1kkq6QBY2
I0kHBHh+/CpFmxlMFwT5/gT9M7fouANbKBuyfubxOnVk3Y7D9fDbvtb5MvOcZkPN3VXJ7zkYDbiF
+WIGn5zifh4W0oW0JWCkvn6MbbaEH/eug3oAzKPTnsCvkR9EwBK15QowITggHJzUbKl5m6Qub6+3
+/V9f5d6+A14TbGkfL03wMCXUxFgHcdoRgu6i7pzHE0Qe1WkiTxMcBHcW+4kJft6CNaBDtGfo3V+
fdG77I+RAnxFoZFNjueXddf+sSpF5KasYUCFCuHUVbKv/XoIXlsvQI9bQcDzj7WtuXyRQxkIqUQk
63IYbMd1j/hwXKFqN8LV+fsVTTM7GBoCUM7BtCinFUiU4vH4fVPFfxrdyMXWufSUrJ5hAdNpKP9Y
Bmp90vWN11bxcLQhsejQRHippIdC/fRBgGBlmibOYsiSqUD5PZvqIrb7Cj4232RpK7p9vJ9vkFDm
RLxT5vQ9FG2zw9LM1ed0YtfNSLhcqjeanygi02k9v2J2o46PVbU+H+dsXsY42uXbRbLM/elg1mub
Ht2HjADcPAYh29OUH7G1jMHkzKO32jNoUkm5E4kabXBLu3lZqfdZ6KQzoarrVFQvTCU3ueUYa7PP
H8qDMFjakZTjPBXCOXz/zhL1kgh5Z+Pefa5xQm2WFLqxgfi4Kw2A596DHA6ylV4Fc/28BO4fPsy9
o9QWfc4k9YaESmkjQKovJP3Rl9jC5hzhtvZXTm7bS+2scVUv/eG8Ai3aiiVeJ8Ar7ahLSRPcYFSb
NO55GClcwoZOW4oSAC5Jbuxozex4dcaoZ+XsclM7OAOdpg2gAOnIbDxT7MfI9dfHHDHTu6kNaRrd
hqqtKcbi+dgcWEFogNa+TeXVpaXNnzNi/GB6zdlfusKvr1AaFK2k0tQgGAPcTbM82OmkLZ4hniAj
8t0I1zeY89MR3vjme1rGGAXyGZl2f+ny53YQ/Wmo6AlLUiZXUF0vA0QCoRgRouRTAulG0ZLP4T8G
s39wvcZtEKXtI0O8wnDQS5I7KlftSjmX/PnI3WdfwVLgAAc6RWuSe+R8WT+xA4iFJt43t2hCPU4G
blZ/++08M8Up3eyFv0oc2iHRDXeQdTLrYVcN3DROjshJ9GmB7V6p/UM4GZ40HhL0+8Mcft16k3MI
zzm727pIFPYykkpKA71IcjwF54lhxH9+GM/6gtp81NJCnUgNcMQmzUNmNlpVqjCk5YkAP1MvxfUc
JPnz+cO0wOV4iZcLAskDnNjdL3FRn0LQVtQ4ej8on24kEKqN6aNCfFQV6rs0rpXSWQwKZMZE2d8A
t81E0Nq0W27YnzJrG2TjwhmVI53iGffNw1Ybkp72EENyPiFcEeoHwXvZ+Xh19sSdJq0M9uMDt9qm
CtTK45aUKEvAmwcY0cwCLngMSDJoAauIQmy1VxyNTAPlVZGZ4zwZe83hc/BMoBfBO/9Nd26WalEB
uiEJKfuQPqbSgHTVwQptx+sqO1fWZai06YNtN2yytHStVO4Oo6fUKlmK5sQojKGi9EckwUurkynq
IQ839XRHebaBfGqQRoj/045LgtbwmdBPw9UcAdNTRAZaK8IngJwnCL8oV3UnZhj9Gn7e0SCTKOa4
UMYKj+VtH9ASjrtak6Mj7cBQ0aNP4ZYT4FeLRBAiGBWN0efTDOXpOKmUfF2dhLs44qxTxTOuSGz9
NaJu/SeFTkEsVBCbq7X6n/+TOCFWRwzeqXJ70Mc8PnvxQ63+0xhOsRiwXDLhdnQlNemknvwgaJQ3
Ai7+Ez8iSdEWsUAXbILtGGX7UPUxBY/zZlZpfm1ikRih4s1+nCLY+/ZtifdB3i7irE/u9uMn/T21
LGTJ5t4sKrvuFmyJ9RP0SYrDudqX9KENvJbTHn4fSnWexDYhiviv0ABK0J/85wkEUFiDfPFVfJau
gAy69cxHv8uLVIcCk+aHaE1TvMZp7PIKMhKkI2p6sHiBSIxvnGCRhUfvPz5TbR88FUh8LtAe5H2z
HVZ+Eb116qIY+1fufe6wGTl0lnJLuM9sOYhY0OjRFFWuUWMY2fV7FDoyya6xsX5SZX+X+WgfJfpD
ZO0tKTE0zri+tp78rfGgmHGiD6JyOM8JcSfnLwy6oQHbwPH5hO+ROSBXHvLrxfcdkRHf/MtQuSic
4peTIfgdGGLZBUn4S2ULVpef5O/zkZIaiD1Ead2VZdykZWWFJR9W/YRFaJTssPis1quRKCqPBuEk
cuPnDWUYMH/Y22mVh8w0ZBsRu0eQN4ykuu0xuJTVTWW6l5A1Icehsq2f+FUMNNqS1Su4LkPv6SCp
Td35w17IGIYP9wQKSFdJZyxY3mbavtTfcIgUZog3yDB2f76FMp0mg9kggFyecBKhE5tYQqiOyc8h
i5yGbcORWheY4SksRIgvruXKgYAIwL6PmginkZke97ZIPwYfuMfl/ts+SCVAOIZeSY20tk3ZHhTC
wt+EQ2tPWQSAuf9iN8ZRmcNgjnJZLqL0Xn09cNHNrTj8UeXGnAFYa9BJwNISeHnWqkNSX2JVbAPi
DUzi9nZjAol4eJzQLMOAJKDC0T92gHDA2ATJmuwjycUJEzwsUFLX5o0fDrrjitR3NMuz2D88CX76
fbDj9wEx1t3RCpLzjc23kuNfh7hKX6MeOGeOjuaeg1SDu4pLrmWxNjBUxPwi6VVeXrdtpjed7WIy
tqHjN5pTg6QQC5wtC/8OSbiLEeg9KllyJaKzObzhQ3zwvZS35C31VNWxBPUc2QQjpl2ypdgNcKA8
x+k6ciMzT6NNj1WyyuztzaI5QNvn0TN6/+2xOxbCf+QOybBrmEhU+ulkw/4tRVyQzzPcT0/S98pK
N/kXRRVL6xGFKozN3XUwlguTT5Aq/q8/UP3wskSX/CGBimOPOTWY6sdmnmwv2eir9KArRvqz75w1
Mlff9Cry/DnPZ909m01hZJqVgsC9qk6Dw+I6LGXEfepYzTq3FDwiy6MpZ+1Imcm79jiu5IxZxVAS
ECXC/G3O0WKQ5CTZsFTUEiYoYXm0mwKddk4ppKahaNlJ5D/n8qea+rIWp/boYp4fv6UDjVr6Fg/d
03G2689taq2P4tSGOLSMkY1uerHzcL24cghIkilE3fAWV/tGKqAo/P1PRa7fMbGTvPvVXWGUsNpB
MsVd+rEDWfMSzQ5WYyICODyW4KcOZXw22NUYDjw17dYLEYXH3bbUX+spYAxuaPOH7zAxmObaorSY
lbQa4ImhMv35/PjVaV7ItsKMB+D4KvZq1cFPKWhlZ3ug9tyYrUbL/UVXpq8MxI0DyIP3LINE0rPc
Lp1kJJavTptjNrnNm6SGF+/RrruvB0G8Da1Ffn60usNQOs5IQLHVKhY+aH9iakbEwfHx9f4YUuf4
Zu3bBtVWpgkAUgMRauNhkkQEf2UZwkmV4S7oUzbrF450cTbPHGNlG7P6fiT9n3vTot1yKQ5COrBn
lvNZR5CxY8xzqurYOXrVCBrAcDt/gKfGrLjUHOfJqXPDTBmMQV/E43edhwn15XlKaHuWRq510Kzu
hQS1W6qPlcQJYMUZXpybKYk81wkczLai6VR71sa205HVR/TdAnvqNQShIwdaYjpocU0s9TAMUqY5
/du6Dg1536jd8OnusNUGw/uNxah1mzBqRbieAvI+vfk+fFGCh1FR4itMhjEWjs0TKKCxTfqhof6M
dzPIeYHXVzr6FyEUm9gYNbashoCYnTksA1cmYcu7mEjxiR+HwTXfh2ur4ntu8fsfm5ycw9Pip+OL
9rXaKmgUcW+ThF+u5fuLg1yUB1MQUbh+BACTyBTlWlLTGwLMNJNDhwLzNos/R5LQYlYgO4mkVfYQ
N8iHMpTXCUOa18JMwYOPj/iy2WZHh3PQbOhG9YF+BJ3sMvg/dpB2w2S2IE/chFs7lGc/mxJLMPpt
Ac49zgAmzzTdAI8iGAf5b0gnUeuMYrxBdh5V/5JqAHYrvkODOwJN4jbcR6wBRfOxw1drmXcFweAy
P10Ew5ZQ1EKfwxYa3xl/9LzrqesI1ACshSVOPXqFvXZI46gUVzWKvnKEm4lyUKtaQungLzSZsv4n
PuF+mM1UMVMDBTypRSILL6xVWg+Ihy17qAlTSmehHc+Sj0o9UsXgsxZ9+wTUVpjapIGjooNZ7Np4
SHYmtLGcnu9RD4zXnSjc4Dr7vojTO1BGcCqnG3gcYrA2auOxWneboGckFnSffO5nKGlJjQWu1WSl
p6hcEFV4YHlu3ZFOzy0XFUaPdeFOwKIkuZbOWf1BfNPr7Q9edsfHI+jITXElf0hmE1TB0kAaOH+O
E3rPiciyVSBQ3ubXRgsZ2zmPMlxV2PTXZKnZNs5xUhxQaPrZ4vID8zkb6uU9Sk09lgcQi7/uAU8M
GO+BnIQHhDwrIoe6XrRS5yP5YNIL/+eZkFzqd+MgiXE2EcD8jtqB/Bexhc4O1rnhNk6VtnP7SMji
S5DHyZWZu8hBNAG9nqLxlHyqDZeCA6VzuS5fL3uoaeP7MGWs9dC/mY4w+YA6e6J6HfEvL2tcEN1X
CV+DaiSqGV4btFVg5QUTmtVyo9E06Z6RY5UHcOvS5k7GtnAOvYfDJCKptjt+N9mnE+bNRwZDqI41
CscncMT43YAOLOcfLwe/ybUXqDDlFyw76rDLYDKmYMe9IZuD22bYJM+JNIf2ReBqTjlz7Fn9yMgw
SYpP88myUg+w9HsTINEXwAdDQxnYzrHU6LzNSZXeOdsJtvu1UXtd9lVKHYI9Q2lz4Oj0cx0pxCWU
mJzvyAnJGq4dAItOjizTCaWLzTKnXGWzDe6rPg6HWLxDp0IEyNLRwzWw/fPGbNn0FsIAvqn7373D
sADgTDZ0MVourD/oeexS6ceGJbxPAC3YPfBkrA0my6cOvIyV/KrIqsNr/Y6dkAMBwftbUQnD/PyM
/KWtM+uGvY+E/F6wXyB0sT1cQXL4u4asAGUw3xKdpzk+Jbdzrw55oSCDBWlO223VZQZsBrfd5+1W
1beqFXXON9M7Qrif/QK4vjI7Wr1KjI20nUmA4rCwvvT5mp4KOpF1Fkguc4+qhLPR5rES9zvEqSkQ
RF5L3iJbTy3Xnb6pzVauKZ2cFf0DNcGZ/tgZsG+/XzbyYq179bmsSf3iqoh6BqKRdT72E2d018x9
FDVfOKQCWURF4IZi7gdUOk25spX47GwBxrDNd4QIwWV/6oD3a3nuTCXrHoRP+Uty0ue9wE394tII
5KR7Qw4TxzChE4o+Ld9UgLUyXBvlTiVNpUmFT/zgw6GG7jSCBybQVF6tFTJ1M4b6eJhqgwDX2RNF
Bxhh1CeV1ZVD7wdgvF7mlf0z4Yhxcam9UYCvnLroY1/u0YHbESkZCNwJHR/qZZCf8QSfquH+4WLD
DPf9WdyHKmeFw/D8UJzm9PJYP6zm8mZRU879Ry2AcxJ6SxuhqGGm/sx+qid0FLZSHV7pwD1E3a4p
xX6nLKbeqp74Oi+7+soTOIujfPVM2qGRc3e/joMqbalEADnnwkYfG+QOPPDd2XzpegIpZqU31PDr
Vwfhoaulc8pEC1waZexLFNn7lVSLNBeaRN8tbKYOAkSamO6zZy2DDtYt07pmbdd6GnXjLxnt5kYI
eAw6n5A+0AB0r8DaSM668Qkfel4nGBeFIOhADKpL9mgFRkgGvqHD4cXJeA00lPP3E4g6FCzdXvyE
gpqqgG4cwhKsWA4RXyQV7ckFOnKMmeA8TFwFZae4AWt9xRCi071AepGFkkWHxA7zs8RlhPiG1rc0
Zks2yOhZvoerzPRPPvtfeScsfFkwC4SJmihDHc99Jo12lEnefNYOgftTB52fWQrPwj2hHo87oHuS
+cgzY7/lsVOoMJ13bUvyhHNwqjeaw53c60ukFmhS6lMU9TpzIlhBeCjImQ+VB4TvmcL3jOtUZ4Sr
j3JGaMSUBX48qONZ2WbcWl5vzoYty4nydLygf6fudK3GcfnQiB+t830BsC5vLzYV4zVdFM2Zymyv
+p6Xp63+Tf1Fl1C9OIXaPAsTNBA1ARANOHool3UzLLJx2SAL261MUNj9YtBPTBBBi8WAoSXmESgM
f4gRFQZIiUUXNQF3NYyHnjs6KqnBugNJYvHgL0yrwI527CcVba+iqXy0hhPXBNqouB173vwiQQ6a
IkPLZ8Zw36T8b5EDZZlfH5wvlrT7enMtktYIcxRHGdJqtofg4vEGWBW3xG4uK4Ckib3MSTb/acK3
w44YG5aD7nij5tjEY7xxFdUC9vcRrZKYBFz46VixH1CEndLkElE3Wf3cu/wN1hQnpxholLBs84wG
VP7sQsiLHMBnijnWduTShDd0CwcovhRvCFr/2I0m7h6RFftei7SEn7EDr+Los16RiqJg2BkuTCzh
r5WNtvMmzk983EVU856O+ygWDxSyx2cSpQ9KGBgMsdUP8r0oq6Ya40jxvZ7lqdfEfyUHL9IY4oVu
Re3Ja0r/HkNV9jAUuPY0G5kZMCGNKTIRceISdH3Uu6eMTBrHo/1CxUWnY6SsVvSjl6mSfZCD/AD6
BkTxMO9wlOQJPPKWHnSKgI2NtI+p69/faoHoeieAkEpk9uFHfdIEKN2ie1gPNZjaILd3ZqWiyYHe
LsPfdmUrvILNq5QCPeCa00VkN/mHY/iJf7QeUNEHJSRjcKBTLgXjsX9N2t75eOElQypxHbbhq12r
hRoNGIwFBD1MjPxECxo1UhPi+cSDBM0zDdStyEc0X3blwKnRwNJwrlNrsSQCsBCabeNbxL3zKQIb
Mz4afLVeI4Sz0drIg4w9PzxYJ+S9haMBF9/KwDYBLuXbSzH1IhKrnYWV5l1lMJS/PvApmWh5VUl0
JCZnWDGTyaOTlopogLgN4tjxmJUPUoZjxizCSi3ZdkTvNGAVzKCR1FOCdKb0XreiH9HI8dJO5yOA
sw/pI4TVXnEMXTkUXvgMZsgTg5GUG8vrMSVBvWW+AIhyYTvFfIN1kS5tr1L3R2gzWyXPOXj+ezwR
U0VRu3zOcGUrMdsqO5g1RHZuVmpDMCiK01o71GaPKNtcnnnHzXewQsUSx0lNe/CG6YaM96Y2/zMV
hjDLIv105i62+qgzKJwodHc0jQqgZhw2sdv2y5QbPE5DWSqdOcTYHH+z07rACTQSvkDzCa/rXqUk
7naIyWlu8Xd4SXP2QEIuiyFnUe+ZBKsa5RcRjR55B5E4CjTzDJIyhDVF9JGxZQeJw5Mqyb8ncmL8
zeL7g18v6AYwMX1BwtL1bVwS81Zzk9PEzo+kfBimTiXfZsE4jdBrqMBKDIm7MznDtZAOKlDswknw
MohWv0FrDmme37IOSKDrlM6pclSAFriiqur5E1+6RLOWNnk9DsutCkLq5dy749UBXsVEky0bIqmZ
N5A4wgqPtyXVQFeDZ9QALXyHufE/3iC5v3zlMCAF/izfzSSQOTRLjtn4w9qN0F+hlrDSnzsThOed
gjXWZ3s62On2stguR01zDCfTln4Z8PPzh5YdWo5j30ES2qdDjZ6atStt8bK3bhz3bqEsOKwPhDUB
xzQIRauBu+/VePzzOzlsDONgAkfwGgb5QDkWbYW8OxhYtohv1oVvO+VSdV73A45JTYp3yLndDKUZ
oGmO2ouEbEP+Nn4XuOfsezDOcMON7NLtX0J/Mb9Avm8B8wA4DlNr5V+xV4EqEZfgGKKfgvNg6liJ
xAn+HXQKqH0PFMAr5eYhIpBgYP1XiPTrvGKtPF/OKcBdGj98Q543Tgxthp0Tp6/fwGX8oSEKwKay
GLSIFcIP3AxRXWIEUhJhJvRxEJSne7/wzKjTuQrWLnMZQs0Nflj2Nb9/b7VAGeX3auTFBsvCePrK
uzi1TGtgQWailvH7gg7l16X35T4mi8j3x9IMuJAFeqRAyrkoZRw/NUZ7X2ylD4TPFEwnsYwHcnPZ
rYWUwvn25UtFWKQlqrgJJvjJ0ROeP+x8EFaeCnePuz79VHLD9V0/ALTG8kz+Lz0D/Ng/sebAwoex
HpXO8ZYPIjcA2CVuv32PBKC0OY2SXstT4yeNftL8Um5ky2maiQVc7tQzSzIwlQ3H4SorfXNwolMD
5g1wG2dPjIqHwRPcHrpvLaHTb3HlOC0zDkYwIuTFoeBnYy2rhdNu8FkQrPNQJz2yD2eq0h8Sy8Fn
OMmS2NICkXznbYm88b9puH08Th+lBeREToJy91MgPS7CoWzioAYO+0TlwgA5Q2LdzFIMiTwHhRrb
aojmXVuclqc5UL1dBihMTxc137PqCl1VooS7Jww3OCYFDpGLPlv/HGGq08EFJCKXr4Ck+O20zbY0
YzLlVF/de+lhQvM0AJwrGn7eCU9InQyxIEiuVzpmeM9TG7UhxUvWQ/iNEfTlvYSvWjrCInnP4QrK
XEfwwsff39fIAnwWDzhNUiw992N24wrWfcteXHCe06VQ8tD1jL6IA+BTOiBzrwngMxaDkCtYy0eK
z6PZP9kWVT3DF6P4ncRXecJI34TdjmeNfbV7FfciqnE8Bw4UMXn2G1xKnjCoCFMlwDeF/J70KBdG
wOPrD1ebt6+YGiPPEPIx7CarqlpqxroRmssYHceg3Gz8IghbcqeXJcklC7scXd2DSaq/wHfs3Zxa
Xx3s9pZAC4t1Z34tKmwo/MxABm1ElXnGmxD2a5mrQJN4UL7jRLbAlxKmbS20bVJPo4/xjf2G9KWS
Nwk+mZdTTWJ3xjj92iGWQg5ci0v0oUIjLFpegClnJ4f72lVmtLmEHRlHydgCwx4dvWeVyCfTc9QV
i2dIY4H4ZyBs4GO7y39rIJbKVuAxESkkms2FvTwmi+pX5XlLPqD1GifuYR3Dm/bWAwrS5Qz7ZruG
dhqU1U+/Drv2I2mNKybrioD/Tkp5491uq9UIoq5AcJ9mIjLnE0pc3VCc1p7znkQcANNyWh435cIG
yX0KbpVEDoqbhRVpuJt/HMp0XhXgm/fcZGL/oEqG3YspYPtOF80qtbNpcxgEivXxtkxSOWsuvxxG
MEuLWWjPyuI1+e69SOTEaVWEnKjE30Y9ZA/AivZP/5grG7DG9kqK7i9mwIc4NrfUV/G9SWHVXcyw
j2AoZdDxHzzutZNRLbBwbzU7VACvT1+fpLfcOLjQL2S7rMdVHjkQBkPzfA+ZxGl8CYywr9WFhH2n
rkaWlzJFVyDCkZyX64crbDIrYwadhAMi3bwGddeb5TU+uyd8DE0MID07/3dQ100m8dqr6tEDe7Ux
mlEoSIfDBNZOM3G07pvdxDV4FL6oVYhy7sC6BgbbuvDRQRgD/wkQSNuDA1weT2wbtyMUKHqjeF9Y
OuSNo6ab4XMHpndatodf94sYPFaUyEcY+f0J+vXV8f4a1BkSz3jZ6FBs9Hce8q5wA05c+IZ/d35F
QPRHPRecoNx87xQ0c3vfOsGgq0MkvvRbO6cCzJ/+zj2UzVYKwReDP6zCESZRdfVyYxfBwO6FlQNv
5IaII9BWvX4ErwkG2NomgshjuYUvi3F/U+W7n5RljPPg6MHk5rm4evzRckdTZXyhxtt3idgQe6iB
ZGLYGwM2N+c/oID4RDQNCXPDevVsNnRxUF0igwG5hZgyAHCjYU+y84NzWuxpL1JCkGOgyMQjssWw
7XhD8CDeR5lmk2JscF33435U7XqHsitGCKYU4RrkBJj+0K/TCQYDeGb99C+zHlVhFv39JST1CNn8
pYPmUNXTlpBY0jXcRuDRhSpJHiDw/QFSWRrVoc8jrBQ+a09Urnftv+lnCLA+bAkeutA/y3WnJMPD
Zbe6Ntic5Bd7u08S9zPrAV+Rb+mVAso6N1lSAmaLWAMxxaA0IAz7y0bp7p3kDQ6W4v7vfj6uVQaJ
FT+/cpd11uLZ3qVmXFXaOYixcm/TgjNUvHVjk5+gZSRTTuGHmsBgNfZm5CsNBik4xb2wE6c2Mecg
Tl5hwRQiBBCCLJe+Dq5N6HTX5Iv1LZyPfRajfr6ghcYob5y6FJjMZ672W7k4p2Wc4KMxxP/2YlUI
y/7wFyvWZP9kfmOgL9c8A3f0OT+f8KW7dKS8EpWorb97jOVxc270W1DBvbDNuujnefXX2YL29/pt
BXsj6IVQwiTSyTEj4fk0+s/XH/b081hSozwOL/Ja/a1AiK+X7O3Nu8os8i5oYjzlBE1ebZS+H6KF
4iyeFmatwfpZ/V4pgwIvSt31UKAVhTrYAc8vqPVXIPHsW9ICKQjhH6Z7+jcMH+MB+kdJFudoOiKJ
EM9s6f5BG+vkJG9vLSFQOQ7X7A25a9nJfR8u+DmVB28I5Sj3IQcHoWFCbsStUoqr32HAIKzo1r9t
THPAEvJz4RYDRY0sBUovLqJgXjdz8IZJyfCD4D9c4i5hlgYdp18YM+ThS/36uYd3W5jr6xLX8EA/
H0OrLYz0RqlKvVRW+tYc2lIl/B1itSNal3yTIqQ6UPeQJvmVcYexgzeoawWlf/eJ2ViUX0hO20Ml
JrTQqvoY12TtbM8NvpPisyfoBS62qUN/blbYgtID+qodVg43BN55AFRp9e669iqL4x35GrQvILl3
t7VEkA1smoAzd7Li88t7txMEYsOAxv1zQiU9r+Wv+zR7iyxAAob4wslcQhF0ROuPEfUeuuXy27hE
rTRvacDmKAnpt3e0xQa8BikWB4EsaD2Y1ElzWe3Dbu1VnS6qXsrhca6ampfkARnCceb5EWYB010S
X+UUjrWdeM1DV74HTfSLcqHgJ0VnH+EOdCPLtlrAqJfW7Do07OKJduGgkDN7O2iuwJcq9M5CxJVE
bCxn9J3HksZnHmpRUM/9nLEnvFLSJQv6Ed+wKyFOoRQgStIc4he9UV9QW+KTReIbTjFwD20Ymy22
2BYRMXoGwDTnox4eI9y8hLP41i3wrGHbxZ2pqIhDekpt9yXbqUacoGGiHR2488zu2qOeq0YvKWWi
KXLus6wEIBnDy9JPoUPzx5Q7D6Fv9tP8gKS+c+KtIJFPfVm0lw7CuKYpCP7sN4whIggYLblu4OT1
AswX9JTBzcZL415RzC2E9k+2ZH6x9KX/O/BZL/+uMasBQJIXfQ/u1Tqd7yICfBhtdcaryI7nKt/Q
i+A5tFwxKiDzW3mMM+unURTaRzT20kgfMe31gKVjkkrXkWuthr0/uyE65TILSSG/fmVOjtlk7Qfr
X2yokA7GTwM+UfuGjNAqK+0RfCTgUxY+a9nfoT5n6QjACqB5hCERLmWp2nur+/Ljupo/uDYQg0ye
NgKIs6d8DE5koSMxMgdyLE6pfrxuZROBN3UFELezwuP6Nj2IemOlEDy842w0fbWMg3IUV8VV6av+
IbMMWRy1WbDX5Z9WdRsq262lOvpijMPEMz2/RQ1Ek4iLhe+avAjc8gnlwCVAhPjxjllmvgNV4BY9
x7/VROGaasvTExQDLj6KB6uXWf90ohc2iq6gba3NfQQ7ZiJA9tAPbBmTlfofdHKKwprVZViWFhQP
S8ufF4EHizQoz3+PfuStsdU5Ka+LQEuJmpw2+rfxK9HRvKyF4IjSHNRQAytqMyAxFKInw1KSqYh+
71D2UwcncKVDtmken6uhvjBHVWEFo2GKq+R/UPWU+UoFxU+W6Yntct9wJh40lML10ZHlfDZLOfQi
Fd/f0Ircij5x2qdJpGSNTdmsrbXknX9bPvK/gVehdg6rxTHBb6ELTbWFr7Co4ILc6b258RP3ajfj
EtMPjWMat8sX5la5OLJDHWY92v4GuRojOc+hW0IBSbE5jQbNc1yuAU9Euppbvk/WzYuxaBvSK3jM
xqTrE3Yh/YRGGBtu1smhmKDufyQw9fKljYWk7RZawzWgjGilP50Wp2bYMsHsSJhcKFFtcFKCoaH/
ENi1eQgvjsOZLsyeW4ijZUKZiaz8s+7oWN4QJMm93m8j8O7gZ6MwsYK23Fc2BdCAf2BYLmKegtdE
QBDY/3kZCIFr/Cl7N7f8r1zyQMRU8Xi58P5Oc47ysSei8L12RNvzOaLQQbFDjF4758Frt0gaRDR9
2WAwD5REcmiRCFNPJ7HtcPer/+ahg8VurMCuWEabYE3SKflqgY06mFC4Bw6GuS2ElF2lFnF9Qik/
1Xs/8mr2sG44DBJCF6wbO1aEPZoQN4cTuVYyQGyIBYXMwOm3sNl3z22Pvotbg1FRTvWZdGpk3J8V
Tvsm6aqLLyJx/a31sKxeywG8pVXBBRIUQ3BxqH0Sp9fWFKl6ss+YPanWjKf1JKkFQ5JDVUkqgGjE
6ko5yLf7SFvIG/qdnUQhQNZuaPi/kYWcgIxcwYaEPszNCUnUyYwSRmxRuYkpQzxm63w9MP7QFOpj
t7Ny7ECJub4t9h+NpxWfsQ1NUQ9jIhRF8hFAgroNJIfimrcbrwDNoqFP88xc18OpRMsDt02UTRWE
22WlnYQQbfxfJW6/t9aHnxKP0GAQyQwy9AsngEMyttXl5wGOR25jFG8BZmH7rRH26s4Vl9VcoKFg
P7dP2KDcSVFWVH/m1N46ZT/vUekvs0cyIPecwrLl7HPxKGZWgQ7PaePO3GhM+oLUOWvhbxXjM3TH
j5LPWawvQjtLTUZtCnPL1u4fpMijoF1pFqSw/LnWiT4Rz6DP5+ULZvP+MmqEFIPJcGunN+QCoB99
o1hS+AUrkkTUlUE+/XYeVIkAKs6Jh0ChV4gkzUDwt6Pp8TOnAb528dwBjkl++vE3AdVGzZdl/pAv
7IIMI++b/L3NYqJ+dwCV8OzEwd48yc66C8SYsq9SrwlQt/+MNpx4ZyX74gIz9OgydLJkrB4+zLHg
yiB669OkX6D8ARglKBchYXYdGPt9KDU1wthtp2ZvOZ/6lWlolVs3zpa3K/qYlFEr+dRRlopsI0n0
eZOC88X0B2jeY2MCD0DpGaLLyu2frK5gZ0N7kdQOjyQv79S4yLfj+uyaRVgnCnXrSsY8PqdcM/9X
o4Ct3MtJmbMurllYWeYaKMhC5duP4K7+eKk7+P6qAobBJuB4UGPZwHIX+QAsSQOFnWNP6AkxJj80
MqcxW5oRSAaaBlK6toXIieAWBV4kasdF+4huMPKSNWBeZimaWk1p450U30APOq7WY+VzPOz7dJCL
0qlLqKzspotoJnZ67XbPkHyveIsoPNLyyPnan9ASxRbJU0qg3QwLwHvPXNlv2th1jDWnBZ5tR5+Y
IogNGJ/c3oKh5Aq29M9K6JMYvHcIdtJA7cvQ1vX6n6iOP72j2FpFVgI4V8R9dPtyYjR6iE/W7qW2
wfn1h+gGwM7OpT5GZPvgwNirT/ylX4NG0nfBvcSxCIOx2Db9wWK49YR6Uj8k4ljXwSyXJ9teLVj2
mIRqcNfUqSRnmmhtpdrwWq+7f1qwp0aW//n4xRhi3xpF/FkDYZC3z/qBNjyyHNgxlVg+Yv0qJMWR
3A54QVjcAcyb5aTXE1meFXbFGSv92JoWF+Xney3ssAo2ANPTJyyZpUPlciVQ3lb7AY5eJRE+5OCj
e/5xA5ORaxeYddV6AfiHXc2uZ4CWMCmfdjRjeObZ1MCDF8ZE/Y95zVmBOefGCmY2Bv+0ohoEoOJa
WP1HHix3SaNoAZqTBrxsEcZmAEQ5hJQ3weMSEu/IqHh50Oho+5g72rAikL67TdwUMLhkN/3uUicN
0b+xKrwqVih6uW3TT2ay/Z/ndEtRpxNxxQd9dSxytHJwfoNYReX9j+DkD9oMpJXzRlJSesDa+ewg
xXImkC5HRedsHyzboASo0nSEuD+Nhg8FfwCCLg0umXZUtoU0Y4Lajy72anPjICsliyMys4whT2ML
zU2HZ7O1fLSt16vpQLOB0FVDutE30Ja2X8599zSE5Hx2xiCHpGGnq+tvpEN8Uro4blRQv13YMP+l
we6Lh7fOny17WEDVdlrVx30sCC27vyztsR/QPGXc0TNEj19/rCCEnam4UymG3kTWvyGUprMwIs40
5h4iLTRsnG+IKAQjvG5NHqDOzC397bvmjWnRXlsHvL37FOibt/StCReABGsCRxSpaBiH+LHWK7eA
M8AXTn14Mm9xTT6Y2j88T3ToceBN0JXWDyjOEJoh/NqgAr5sfJVeJDDhTmV6CXTLOdhRtyYUxy9O
KZRvxe9JGvkN/XfIVrem54uN6QMo7G5Q3l5kAF1P/yOzhnKSg2HzUvOdVtg5WXggLtHT99NlUqK7
Yp+AD0kYSqB5HmrdlSXw9efjvOJjuXWeT0PnKR6I2mvdjf2MOLD+b4nQSx5KP49K8ZRKZNQoUZOs
Kr4rmC4ludJgtpuB+U3IUgo8DBDOrs7Gjmr2I3e8/e0yF+uXzyP0SefRdgCAiqm3MaeRqINLcheb
7OoztwR4qIny+uiTPpQmcGqP9b11eLTyEFfgPJSNom881Cmfuj7eUXXvFLWzJVp4/Xxy82601zyV
yu5zqFZTEPDPS9MpLaz4Oh0bAMSNakqI7Rn2/qkKDxjJHg6XYfWxX0xSFJGczWopucuWk+jPRQRn
DKbMgd9yPx85yxtKXp9+ranz82XUwQiJ7uxC6YJ05gPGDqnuI75FMVVuYS3/zGV6rcfdx67jcK3k
nA24LosYEBwFy3m1yleGKteLnqzIOQmMDy9IN0AcKnVZj4Vvzt/5d4V0uTnulvxnp9OUfL9Fxwel
JgJ5FvaY+Rq9Fkg5rESKh2UWZ2lQ7UM+A55tuyhDjltZVyqu50reX0prdBuBMWesWOyRZ8YPVQgg
I8f0XZAdofAtkH+z1+uxCFNV8eh3+ktVz+SFA+whduLbkZPvz4ySxh4ecTC+E83YZvk8UwvNgvJt
zSzjj4vv0ODNLkiOlsJBVlXoXchaoxno6HP+w21A1m4KoMnD3/EQ2+cQVvi0P858VjOLHVfNLOd1
OI8cMKDEqaI2Q0HJX1fAyWOVg/c+ItuvpaXueibelZA51Yc+8qVukNtNtTN/r/x8Ps1zfW8Bq3xG
vMn/MDOuJm/AxmVUzazYsAQoZTfph8ex7c6bCbqPoRj5VW+WSrnbyU94+o0Pr5J8PT+pAS+Xt6Xp
pGE5Uk37mFNgQMbLCs7jtmjZxdB5tT9RuJxHuceJq1VQifFtdmxmfidM8GLo6mQXeEFYLzLIFkAe
VLdxJrFCxUDkwBDeafgwpQsTLWnugAGfhrpNdXYJEyJ8iUIrDknHWhfXbq68Uug4saj8dYKTDk2t
wxT5YcFxLsTzRV11pQblYmfJspGzJ4FgupinNS8aNcDur2S7jU/yo++9iVDR58I6DjFaLndHqbEX
Wr6pHAV9cK4PXnfvYvkt6psCmzOf0YuXqfjF9WCNIAhHwnf9odElqi8vDgnZTdVeoMAG8cx5SfXX
YqD50SOUvKme9zVd8SCKJg3s5JhlXB954mBxywbYFzT3oaJq+qdJwToOrsi3S0ogFW1rZ57pEpXJ
WvcK2EHg/fXve747LQzkw8AZ4LsCihcLGEGGBV3hTU9LpV2iQWPoE/eb+bkcpwm1daPDvN0ebCzI
KUZKLCLDpljUCWVHUhv0da4AVydjQlKoZrCG7aVnvl+iDfyutwZAk8bBG2FDma1KlQYXoH5HeDVY
BPYzdMVCeikmLe8z/cUAV1aKq8GYq+8nVJwZaEODS1A+p+SPVVvMBOehp/79Ij4+bFYtSkCXd0/r
jfp+hVn30HMUW7xnd6WHdztbjl8GQruV6D1SH/sQgwaVGKjX1fO4jl8QuVXSJwwhHj4JH4CI3BgR
XXrmWg693O3OixfYCWMzvd4ABPZUubntce4jf3rkOSpkjiMF6d2tVVm/T5ELDU4H1wZ6nnXXvuLc
Lf97Ah6TwCrmyQ8doxMDOY1PGvnyzVcKMMe6CqErYHADzGsA4qWDOFwhTDPZRp8nDymWr0IJq8Wu
V9Sgq8VZzhX3rzyubUonxYEMosWCk4yLZVIAX6lvnWrfqXpj10TbOB4VEYCJhwgClxyQvTQ/zv//
GK9/Ro7hEtPfgrCpECZXsc9x6jckK3s8g/Sn7JeTyWrjINk7X7fOyWYi1jihFyZzbfg4drnzVq4g
31Q2lmVEeSHPUQ7/YMM/86db05weHzesdLRweZCNxvyg45PwIt62fHLCdES0OPchNcyjCVfFVo6b
rpDZ+DKsXi4XNVpF+MuZjqeAgPoan2E6sPJaaYXff0iqohKoOom5Ii0lbDSBZ5Tbx2U85dS8AKHg
a5GnTtExmtu7yC1OHyDwuDsnpuAuJUWVkyYWygIvbIozgp83948YVnlKRJGYJzaY1WyY7ej0z8p+
JvnGejmnB6uhSxJ74L/soDrtjl3fbmB6622iiGWJTZk2V0Kt4jX1cPtL8xfBuTbQJ0LcabDEgzeU
n1OIB1GOeJgKXaFy40AZ+gRuOBSpjDJ2CkKlZmIJPQ0ZbR2XfSVp9FZ4B8tndFoi9Y6p9Zqz5bS9
wX7HZovN1NLLQ40e2YBKblOKKTWwhyjJsKE3Wdwl9BerTVRzwTxMPO02PChNIDck00kdZiEOd+Ht
r8W47KNNKypgH4h7QcoGVjRlZyD/FHok80upm9oI/1rdRjfHWSHqOeOBxly9lrFwjzzPqjXGk4e4
vVtQ7Y+g3SYjIP/Tk4Xo8DI5aSK42WHdw8aAYcHFUSk9lq2RXE6yDLafZqy3y3yFOL6G1uC6BxdZ
iTjxMHDOPjSZzepS0JMDUTo3qh70buj0mAEy6LD3ecHwk7d+zb9ELmY2/Fzm1/85tGffHsxV+ulv
Gc3LeP/KJweh92DQKR9NHqAFow1rghXfTErr45tuPZ/FIXOgXsOoJ2w8NU4ogkv9J1DOTw3Hx/BC
bXtvhLSzhq08gIoaPURLShxUm4HPqQ22a8qFEGM25vxlFqVMMC5kYNKysecKcvymTWkzC/baReSX
kKHP5MASxBrGUbS+2psUi8WlEbswc91+SSFO4ifOzPYCuToFRvgIt1CCJ/8a3K0SCvC+Xwb+1r/S
ZlN3FollftLO7bvTrdEStOfkq97BfnYHISSP7w4IEK8vQOyfOESmYQTfBC1w8AGF2ZHDoLN7MaTp
GtaMntQqRDDZG624ojaUawamRTIwgvjee+lVCYju3xFk5eIusekK6OH1jzEuG8o+BMBax+MQ7MbM
lIrYMlzg6bwpzxiKV1VFuRkZnGez5I8PpLcqXc+6AYHnR0EgyGmpC5Q1cbRO3aj2lw3TYeFn3U89
IAy7Nei/NObq0qipmqLTBm4iCFut/dwMbG9f+BwZesui1xNyvfyEyE0eq1MYXEg1YZTr9OPCHXGG
IiNBnAyzh5eJUEWrxc9rG7mk+jclBX8TRDXAfzmP6KFw2CtLVU6mUAzDHZh+9EvCzwqvHxRhKB1R
uV/mcfEp67i1niwZ0oTgYK5lWzh7hKD8mlr+L645V3ROOdRCRxQXQONETOoq4nwIkK6WelS4kWNn
3+v7TXPOrN6mc6JUNkSb+o4mS+IzNrHP/5iIzat5OsnvX5U6MwqTB/etnvEzRW0VMebbUuT5Az1b
9nqFi1+5VpJLDUPi9luiLU0PEAL+6l+6QNUIVLUOEQBzi1TNUIF2l7arDaNTd1Sxcpe0iCX5K9ae
zqBDpOij49uBdNL5CWPjCmJFGqnqxEkECOcUnMdbqCMyeQNPrCYEV9DhzvTuNLv1tsg4RDnhyKgn
WqZHt+1ofYCvnrb2rxvnqEj/IVs9dy+H25QZr856e6eVPO00OBtJV22g3vBjtARDYyzyhEgCGwl9
7xgnRZLPyNUuSQFNVs6ulAODeumDm0XQNtWiVz07iXJ0IxDdUCwoshwuAWObFcdsxBhOg9ypp2Ll
Y05/lhxgip/SABd3va5Hi8QDrqMe4vUOi8sm4dhIopDGnOc9NtA/XMUJ83H6PcslkCbzJnvE/iLC
QGHWyctrW4x7TY35t2t/WHBb5pzzw1coLjUeSmHt5e5jk8SZ2qiUb+C4GxVemi0v5L2tXvOH97R3
c2iqB+8QaBTUkxaDrktQvu/rrPbCfF+lQ9EZ+pm9mxiYGO0dh2w5NXJc21ww8O4JUl6o0GMIz2yS
I74VTPb6niOBR6w2x5fvPRT9eYfQiJ0euHN5spTT6oPbHbpUOGvGapUtjuZBwStvxoIubRQTFtB0
niSIy0ovf+oSlskiMMcJ4EIxaVYszzqIJsA85L1ruarV+Wax5+GTVcEBGTsr0DFU2zS/lPy4R/kc
ILjZAgX/cADKM6KPYJ2kpKjSZI2PFBjT9x3l/tSkSKuJg15WFKdXIt3B/wL6LGglkVvPfJoc9qG1
GAL/qIm5lMZJcsK2r8IXA0xLcB9wuSMsf3p1R/qmbnijnjDjd1xJBTRU3WC8VMq7eWqB3m2VNhPw
hNrC05ttooC2Nnt91DXEpN61yoN7L1JCeTj9myjy2xdWI0pbqbRvHpx1NR7ru8k8VLmMTELMH9xk
JTB+UvJB8BOStv2TbVmlZOJfLbAx55W87i7KLOBvJfF6YW1U1aDg5b/5rG85H35AdnWx83QWekFM
IBXA1Zx0Ler4e80qmGuV5oKTSwE6IiNRVVY1dRLGtKwtx6eMOZypAnX6EhyPWKZmiS6fUFopzYdX
uoTKBpXfc/gl6zHkgvSMiDxD+VZZdHKSPI8HnU4Ckfm/l/GXp+aaabgMF3qFDiAljBr5rmxAd/b9
KFuexNRhaeSfpIvWQIz4WMDRuU6jhxCaM6htXjdZP4baOgDg8yylDUFEaBQxWQxjdjO1IytwipSc
iOVeX8vz8LvZiaUUBabaxjElLvIKwn3N+XFehblaHiiPgu32APq3ctnhkz1acIENJa5attBABXxA
FPMGjXlRSNFE8HOcEcoiA8LKZsjM2nx7IKvQbyPNA8VWkWel8UgQNdGWezQfFXzJpC+xavhVJpLD
LfxAmTWWPuMnpNBGV+jEOOtxy6YqZ+UyU7gqBZg4Ek59Ael31HTm+gfvsEAhA4VK3Y+PuVQKOrHK
IIcIxh7CSt+mgzJNl4gQWUgSOlyI7xB6w8QmDAM9XHXwcNhPwWolgSVnwfIorZ4m4u/m61+v6nUi
Zm1mV7vhLwhcnnjYQCplqRkfAYCyhFgXFsDXdMH7WsZamVx7jxbPqH7nd0LwFIVgEvVBpNwPfQlt
DVMqgS/Keu7VUCiyLpBRDAHGRjJiW4IvVbMil44QSdrSMatPPtEsm37A01gFDD57jTiWWCrQ3uWU
Vq5KuGpioN2jBS+/VmOK2UMr2OT8IrKKPCufA15hsX4gR7ijLdKhYZ28rjRqkLXjz480MAH4JzeE
rmZJkaKPQWo1iLKjZ76FMEFx3/jbLNVKLJZnEk0jGWSOfXYXJS6r5sTcQKr8U0VELyMxwDk+mHTg
lYFh/ypaCQEQW7bZ05jsyPJIRmghJp4De7EPHu+WPjG0z8iA8jpJygpGw+GcpgfmRGVYwYMYkYJl
ZDXfKhl/Q8kjnx4Tf1aaJl6HRpiPuZmHvwPxei6LDe2HDV3rv4TFkoMbFHVpIZbZl43DyzS+M4sJ
HC3DFK9KRBKesgUIPweU3Yss+FYFeJyB/ZXCby4/C66fRQIYcGEUOCehVZRz3t6ELak+mAu2o9Y1
QQNzLGSBlA1AwEbcizOjMJ/D/rsFjwrxG+11AfSuIS+AabRHc395xysHqmJ0kLjwXWDXsIQzQdQq
hpvty+jTUlu3diu12mwM5Q4JMUn2TblbURYi9wBm9lX5RS/xu5Kw0Rd/vASoGtHa+b6u/pbjLSLK
kSzQJh/5/dz8yBCIVmPtc9Iw8e9Ph+WzG6A17DfwLIVaeO8zBrXFFjUSN25ci+FMOUQy/NtHOdOd
88xcaVPDkpmfT2dSfgjz/cTpFnXA13iu9lIJO29bb4+yYoFlecFvbYYtesrNeZ5HUxszQG7716cv
n8Z4+XlmuXNPnxLPfnGGRu8CD7+cREqzVYJyclFtOj/r2+0lxdUi6DF0ADwVi2ol/EMgi2l08soD
Ve8+2HcSL60fRfyj7MJu3UV9NsoTaTFP4b6IohrSOVBa1BICcArAUIfV44rS8kmqayPpbTz1z/Xu
8sayNamh/L7tQeVj6RtMC/VbQZoMwCOqGzaprEHSvKtvhoBD9LWapI2Y0EHXaB8heK9YythinWxu
yPqvh+yRiQBTIZYatuGEsHPjtTUfQ8qbx9dzM+xCh9dBJU+LJ3O5Hh2h3RAZO2kvTmINI58q7rYT
totdqIAdzzztOIX9ECs6/x6zz/Myn8+S4nXd6YhvCNKTUvW4lQRsrnbu8JACxp7doA/5rxbBd0WP
5FoyITFeTRO9Ro2vmSaCchi78Hmz2+09PZi3ZgJqqIbp/ktjCDmotm+IoY7vRno3D/dpIPJT/6Zm
SsAkANEflDhoP2cX8IenWB+ZMFbsC8efjj2SpgVtE0LPXhiHfOWQGH4MjSTeo+JUBel5MdEqUDLQ
jYBka6M2nVUtUaPKTRNC7ECpDP6qCjEKGlXRmg7t+ajdxHiRND7W2t9KRPgLX5rR1g7+G29p1yk1
iHpGQtI0ALUFx+35XsBNy4lV/+bN71eToiznPr9vJy+ytIpqJY1I36Sr651OE1gIsiYZij9Hqc9s
XEsJaAuU8aqr3AZk9PNYxUOQEwSGw9zoKbvk821/gzqxTtRYqmL84HESKiL3DA3IY9kXFsUn4uJu
H8VgG9Cdw7pjTQxPVKvmeJ19Vlh/wIIoh0F/5ghOCt8ZgsItg9l8gbLGCAF/3YhC0uylmGdz0jxz
mj1cmXY8Bs0PI2TdjoYV9TfbvK0Xwux8tHNC6XAf7m7tMV1VMFR2WMRLB8PlQhOyIVn11krte07h
7C2MJUgJN6hfpGm4JW8glkNQEGymqYmqGNDghtlJsFUUexu48NDQsC67PmcHvZh0pNsp1Yjc06dD
R7fsG3/ONw24mt5C7ukoTDXCxZMNsfzHOZESlmRpU6XX40y1nW24s/0RPPXIDAqxh47R8srOuK2G
rijxGvo81fHxT7VjjKvh5yVkHJ+M1rSm1rufMcmoKsBaYtlPiFIljnWVr/osxBEhU+eXBSHKOdx5
eBBbLTZeUzxe2YZDqwDx46YwDXiZqayb0t1XH/XqV9ibPSKNSBjGiSfTlLUOYBh1z3Vkqi6eNQdL
DUPiVBYJQaSgO+fVd0AkwCQgaPRYkD7c6CBa8nSEtYTjUfr3+BvJp16hh76eml0a0VfhI4SsemV+
sGhtsUcSniYCI5e8vj2r8y/JCLlsLR11K/oBh8mN43jAtJHsne0HzuNOPPu9mqupn2HRaHg7HLFj
Lp42iTz/f7sZRIWocbzX/PK9Rh566eNlqHIMxVpuGvNfjdwSnMu9G3OVJ0L/509nHfuythnBAZWO
PrkyQTSMEiZ97ybjdCBEtX7UA4EBh3p9NOQlM9UqiJCJD2prEUC9ZTOa5iK8jbHO0pu52HTR2g2c
z378VIgVhAt1oUTZ9AmDnwijd0TZJ+K7tmI9RwiafEdQV8yl2LJYzz/X9S1gRzd8lFCRNcVGfkJb
ZDDjqUQKvgv/1Wt3U1ZhNbWRtjXk5K8pKMi6HzoHx7+X9RQBp/pqVMG0IEmYZ5C3uIxsrJMteQDx
IZbJmSyMgxOG+D2uLPhrs4KdFgtY4EsbOxAYkKW4pIp1zncASpKkr2gr0K8xSX+tpG5Y9nYnRYlE
Hb4Cbdd7ePKnWXGe4j96cCYmQ8RlAItgXgPGtW6B76GfbD/ZFgdfHCc5kTE3zlgT8yLzuHadAtfN
dwW8gn9z5Cro9YrTyhtRDFwDD/DMbbuptQbB1pFVvizAH2f5Hhrst8JWrbVdYjKmGz+15DPk9/yE
7KBrDmCLFmNMJ2Xd1D2MS10+iegkiDad5hqIcaYDG7w30J+8uD5wFCJr3MFricpWENSJI3kauHUK
M5a+HwM5YY1TBQI6y2KJu5HMpO7IBt83xmyLMFsqPjO5VWqhzwHU5K9XHMHl5N90u6Lpk2GMZS+q
NhktVv5uAzuPTJscjkuLZ9ZgzZ+YRFSm7Avp+qcRgH25SDfXLIktuRKGIOU8Cq/H6Nrc83KRBUhc
mLiJ73/4/2A+U05pVKyPs/hGlBEaQpnu1qhQKDok6Ya225TZVW8olykfvtqHNpppAnJMIjnpdX//
BLKVb/fR9BRVoAkWGGS1Z8nlszhyTuQ5Lw0Xwxj0QUH9HrHAfmkyzsSRRpcLpz3xqgubu0oaIXuK
6Dqfwb/hK9va9AlosC3EnM66zj/4u53G1mq8R5GxrGO1qNolNqtdAAmcQsDKFmzp3q/Ke9qnRtwO
iah7BUn1TnjaPGu0izRpuF8LEKXFfSMgx+GcN2PiycPMieGZdXIj4ogxMSvuDPGe3It6mlGxeLUI
IbErYgRwiVpAGqpLE7ic5FEKafVcJKK6mc72rpaDttP8AQMSREWCQz1dkBK6U5o2bokRgC6DTz55
vKW9sGneh7nHwXq2r79ZjC9RZwKu9NSN/bx/KDegnhzViYKik9KzpTxqM5qmcPCJlb1DY532TADl
5PVXT8AyU1odN6x5cx+FZh+19OP0dbVtyighiwa29/qxGjFO6mviWygWPQpP43qzurRawIN7CHMH
FxQ1Yppvv18tzNJ0YmAJ8GgUSPR8e3iWazF0ftyEwuJujnoMB3rYOnExvb/LXMTcw+vJYVCxk73y
4uRMOZsT/GtmEI271npPiRxhwUp9F3XFZH+mPs+cey2gMAWwQCWMl/Jl1y8LxyPMNu1gOTTDbAYm
c4wfFoCtjf9tW6MgAOS33ttGs8pvlPiZluICproy9jU9VxF/ukAiJ6hA9Q+iFkK3qLgUV7/ykOSQ
GgFp/0IBfionclD8whESm/VRzMjan2/tllpqsL/ulxn984FgRvJ8ngH7vQUUV6Y8GNmd8lu1E5vF
gY/uvtpS24lhKfNEQl14kC8TRqNAuf2putfIXutPEVdcStKP95kkaptJtAghmUruf615Od0CRaz/
PPe9Zc4V6mOOHuObeQgGW/3d8C4j882ks7kQ5xixz45lyfh28FtbmN9VMT1VHLUuDrdRG2N0Fdd7
Bcvx6lQ/VaiH7MXgWp7Fpti68QnaHiPCadwcr+NmmZ4457nh5TWF2W9W1m6TRa+jfqdHYvxS+G1H
c7V5yVmCz40n553+E3PKIvdNMKCXsIAtF3l+AimXjT0OzKBSOvlQMTwpbV4wF/eV51irHX4qeemn
yFJODzamfu4nn9XjnpYJBdAkPkRryOn4GyCTZxNwm6I70bZH0N8yzRPeh+KJlEOYctJjUbpJlRbv
Fmtwp1GwKJBSysXOUbd+M58lCg3FGXMYU5Ewzd8xIxSk95ptmkB8xzWLITspln5qD9s53MIc9HHx
WKPLZ/4cq/facT5QRhnJ46WYOwyRZehuHHM1XRxzJMcFE2O3N3QZjkTS3PaYmTfvt7oMOktXrRvU
W5+3j765dCJUg871xTo6UR2KVdmkwbRJuP460FknPado5v5q7jW22VOH2wdqLJ9UFK94+5iD+Kva
dBCVnG0IB7nZjshXBple7i8eWg1btzTrZ0M9lJbvjNnFgbb8PwF6GM8HHKOwBSTCtYoJja3u9Etk
/aV+jW6zhiIOrQXf6Z4s9N2H7gSIO8ipAxIXx+8UR6nYAc1NT4AKHUm9GC5F7IteayX+wKGqEDfN
dif50lDPfDKE0lJONfoXcYOzx0Bw6/bKIeg643hR2iDEDc5p1BQft5bYEpqGh61OnX5a23UCHoX/
ON/jiV4GiiIBzY3RSnH5sEg1HL/X9qxuxsdOYibjjAvEPEtG1zwMq/V3iop2VJodQmWK+Ki7dVzm
pxMoPMQVH/ZF+lJG7deMhHmWXEL8Y8S4T/zUapg22qD2bLW6bU1VPWgjxw+++LkgpzbtCH15vuGW
u5j+fbn46SaMWeNgBxWjN/CxjZ57tb8uIu2scN7jKbIfWVsVZZXwsxghIkwhZHJuKOL0P1w+FUvU
NVPCivQWhjpmEAt9XwcjbF6XBxfOwWr7eXDvf3nsnQyUw80l5fZMxPW9JTQ3yfFl4i2vIAsrb+kn
+NxcrL0FsyDmnZjTvYBqUt0DG5qvncFvVeY2X+bgXSDkSAVQdrwzGe+ZKd28LirFipTOtNs8cR1K
0y1Jbi8iuAeSFOuYEZgajG4YYDMoxxYo6QB43m/yfBYcJKCgqwe3cTiwRkZK7heFDNb1nrg8rMs+
7G0/GNRoLyji8Q9JKYkoe0Vz/zRfKGRacGrGQg4Ot/+nDhWTEKfAq+O93t41eT7eGiMccbGa3+pZ
3/j6CDzc1SHhMTYCeAJz3CMod2Euia3WvR+QQFfaWJjIe1nWlovCTtLL8cWfUkjDUarofceRW0Kt
H6xZ6PnkUS+M+OIfSRml+7lTf+YqqBS8LMFYmz8pdaRNkEJddlpkib5V5Iznw7e2eLK19m+baXhR
d8sSpgeeTFSnyLY/m1eyvb2Dv37dkn1pEHxnYbFVySSQDt3uWAL3dZJdpimB01wDfs1N8UexTD22
wYSHYGuA1m/Q3jjTldwHRIz0sZ/WPUXRjhgzlYZYpxVhWeoaCS9xqvGM9l5X8Mqh7WOuycT34jEK
45vF6SiTr1z6mgKYAiTZH4o7Fnv6dqfe7XIIqAjkjgrD6CPDLC0I6VyFLgcvgPNjQHsDnyq6rFUV
yBkQfYlfW4cgYx5jybcWyHrXEycHs6yqOnLhHcE7Zr1ck5Esk9GrzCbsy1mPNRCon2tCR2KKrRT7
eo/VseXIGb3h8PZb5BhVNNcUGJ0vTtiL8QiYKkN43ZuarmDY+rEUTYLOaasUMv6/NWW/qIGuqLii
8eZWLY5+DMOFVg6rXwW0kdoqNFnntF9UWYwz8IdEOcKXHlrw/MSc/MqMTjwZEBS/Laxkaop3Ljfj
KQIfAD/ZFWL79uSPj2LR1DoIWjx9n5LCLxywIs2e0ufrYRBQPpQEfj8U6ftQbn5shwTs/z/Ibngt
Z6JFiAm8cWCz5drEM0CeG5kmjndNxlajrT6MqU3I2+bfvIpkOFXcr0MPq7oiOKnlMpd9FVQ1xP0G
TWU9JuK+1ri3Fdmrq4mv3MmuSLEVL/BSNwrK1i2BhFelRYSVdpOuE33UGlujh1z4bKuEaD434HKR
vZ+0Db6Fsesytwc1K7PJaVDVm+LvMJ5P0NB3UAepJ7mL2y4sewlGwnYQ7HlzdNwf7QS9SEVQhnai
b1aCNBLPAVn5RpxUdl+P+baV/9bDV9ObI97z1UJMKBoV2qTxwALWl0CMYGtO6QRjsFLDAKp0Pouo
Uk2c+WUjuHsoSlzuZzETdaeWfhmUbI3PgMEasNWlu/Oj+4kgtJA3fEGKa0N6Cjk6V05azbD1i6RI
vbrmsG7y6JgoY2MBhTHEvt7XCgj+HLZtO8KcyJpMudgYq+hQbiefJoVmfc0vgCa8KdwsgpCNlI1e
tIqEHhaWTthmXnlmEIDF9D/nbmy0JvG+BBYfkUkQE13tdDB6h4t79gzuLnqh4H1Ce6DZl4eW1XN2
F/4sQ1vGtce2cJM7euMUfSREM/XAfJAy988H1kRqBr95oi1Q7mvRNq0Kmom76VaK5bIAZRovnvhI
AlwZ8FoXQdaOzVjyEp4dT+NwJgw7v4WfMnQUbhHBguFxHLbF2QZJoJwuisfE+W0CcwUAKpoKy+u1
94ARH5ByIXEoAkB3ip7Ps0Yg+9XFXvU63lee+6Y6834f+bY9NtW/4XeNSgvmY5byDS8aWVu08YC+
moIjDdf6cdXV+kt6tTtvJJy3MuyQqPKrzfF2VLJAVz/yAvHAdqbz1XtNEmfNisE2Psx8pIGZP7tf
7kEUIqHJPnyezWp48aK421t/w0nplp8182/N0HtAKDAGuN1mbtEm0loKKLRBM+oqZr4eBrA4qt/Y
4OyNszk7Y0j7hlxFjt91Otx4IeYBWZanRgGKJJLEG1Unx4So8HosQI8Dsg+zLwBrITHakcP7wJcN
AuDnnfAKYG2UNHphiYTH4WYS+MF9Nah3GVHrxd3Y2wYp3wHgtnd4I7xwpFBd0TY2MBUoX8wOl9Gn
YYFtY56NTX4AzHfqe4yWFzrOk0J/eqia5qejv7xSewyg8NQk9K7OkIhpXEe8gEZw9+39r1/ZvpBU
b5JRw7N4iZ2yHai+iVUqKa4+8vr3SxR5p56gF/IDKzgae89ImM6BN7K5NMi5LamwK5xDD6sRjJFV
tUE0gC3o0JHCFFfNHjW2uq/D1Oyly2i7sZos4fhLjXTihI/9naZQQcRqaWrrBrG2o0WnSA1rEVFz
IcKVBMSXzgbRoyaNr4fDJv2hhFhQtBmZX3EPgmhoFkR3BUIAmOQdo1T0K7Tf/f9cgrVv36tWRyCq
1EgJkdIJK+TZJhWilgh+I7pd3NUN+HrH1BKwnUeOxtYnFYN4PxDJw7LUBUBnsNlEdrvwlLjcDsSt
37qWG/9YRs4B0DZqVU9M4Uvxr70VcowSVJ+XmiypU1YlljJ9Pc1mEezkLQKivtJQ31jbO9qnr0X2
YmzYDCRW2nxgxo9CHjNh7B9I721xJtYb+L9A7DWsdHEPxCgML7BS0cTXdmyGZ02NjLJl1UVqoVJ+
kw3sq7eRPBRFNm5HelB2VF/OLV/H86CJs+rfm03e4X9DX5mQLbGq4fgo64Pz0QwoQbfCCIlVx78w
apoide8F0RWOOihZ+iP52o1TljkTBlNvzupnvXAzp0nAkaqe19wg0+VjpF/+MRAnYMFmCEXYqDsC
jcp7x+EUqUhaQUzuFZkqAIb4MFVF5FLhK/efAcspbPBbplWriqZOl6DIrfM6CzsNTvUQpyV1mmER
jvxbUWJnyCO4PVfUbreZnLAH3KM6EUQTAWOZLUBK7j+O3ENcoPanVk8AVpQE95uyn3qgwXeBnXjt
KD218LsQVZWVJBZ79WLpGI9W1YmSDpWDpsuOFVPBgCVrjIFAm6enBmPiilylMK1Go4SN1K7O3NRz
KGg3HMTT+5yPFY7cnUf04wSTn6XqiZ15HPcK3Kabkygy8bmoISA4B5OOHKMeGcE8BA+ikxdp3U0F
nIqmeDYVsEb9PTVlXXDoTArsI6ll7Tr026zXh9J4+Z4cN5dVH+MUM/C4Qj7KT+VlII/4ycpOPciD
lpzM1YwYFR43zKZoLe4WbBwliJb1HwBQ4fwihvDfVVzvaV5JwY2rakTQtiDFCRpl8qIXWshYPRwm
7nAK2Ev2ZAxp58MfjvsaYV1yzVePorD3akS6UcLKM3gSXPhbVKF6o3ZiP9bfcv/xg2PYHDshyIVA
TpVVixxtnRKVhn2xcGk+DhaDevFJoz6HSPH1xXfcYQzVTbHsaKCiTK38E8OHiLXsOsL8nOGV1/Lw
TWpjXDmHNM87S1sdShZa9EaZXYNgLKO5cv6AqQTKEqV3CU99BNOs/cy6ij4JLzEPECvNvWJ/Mc6y
JNMr+D+UyN4Xnbw43OhzaSDhHt2XtQRZNwivTEHptHekxgQw2YAFLNr6le8RbLG1gEpDi2BNOgdp
NEI9HAGRBd5zqhdqEkAzX72IpIpNzzR0tCcuRZmru0ydbDxkRWkDPIPVcksMNf2FC93JmPas7rhs
/f6ji4X/s/bR7UC4Cisg8qejOVajtDtt8vOC1pZQIbsmi8P4P47uhdyrTpta4eOXeNnI66Ah589s
BJv8zUEPgfNtKVXfyLDu9zugWiLJYsdhVzBg+FR/Ym5snK+NyQMeYCu4LTWb4m6aSzXN1wEQ/LEZ
AvH3nOI9rq68XbjI7NBplti9bHIWcA7/N1IhA3KVzNdxcmK4MSju+/o3MObUsNy/7DtgxegSYtDC
2xfDbrxLsTf2rgo8KgLW7nspf5+2lz6fLTO+oN5oV9aaAj/SbKNs6rzdQW3qe+/viotj9uyHhKd5
VN7hNYbfb1FElHYn5qD95LE+ToRaaqtCqkB/ScW7OfMS4fXDWXap8u74q7BKkAhdDUFIrvW6NSXC
GaiN7RBxcWw0ZdQgYgtM4rHB8nNccdaaBkz45P5x7C4EK+HqjzfpFVAUIR7gcQ8p0kPn83a1Qxqb
8Gj5L6vdUnaDQI6BO/fcEtSmNMUH3vnAmHjSNZ6llh01/0c7R9ALIX4u8RinyJJWWNwRGhra4+Sp
rLozeyDyWPUAKgtty7ZhP44bDIEUTP4DBQMGlh52JeDnhrm/ESr9nv1re4kzg6oziFJgVNNJlRcb
YwQhhgbGVXqsOHlwOiWSN76tfsUYIgF/Gh2ymG/5eW6sBvDSu8CE2pc+y733Es/pdo38c4mk+Any
hJsm0AT9BJVSOfD3BaHo3G4bcpcOen8hcBktOgX1+8YglKJzGiIL2ylTYBcYQUDEsVIfyn1GhcgD
EbbnZuCjLnT5U2ofqn1ItP05s7eS9ETjCwRAcH1Y+P+Af9x23lVu8cU9nK9N7ABwrAY7bDGv03d5
I90ihxY72kdvKsXPstm7vrEA3XzoaEPLcY6yhaIXd+9hzCljELj83bU1lSrDVuF105QexcwkDM26
B5WvBsl54G3U8J4vJ1rjyl7uwAJ0ojbdb7hOWLrw1z9QfGipTAiPvxJM6jNI/cymVhRIS0AJAXkc
ClTWxQQEVIAttIBkt1iuoaPimCHJ3CqAJXyo6lqoFlQEbjuwVq7JXX3BhGEcebnsiqVQnG6ysGAL
pTsWT6wahbB2U4RcHNEnXwZzPETy3mSVLcEYm5q/V8MZORgjrX27mKOP/ytdSDkMJ2BBohN4DaGx
52OUKKGosqpNPNRJ2RbrNoc+BchGdGiJF/bTcGIvwlM0zCMTXzlFf1A2xKa+kdauGjPjmxAD/seB
SOFoQfGTy4DUe/FWe4BgJd2njOQ0mRTBiTT+IvuBvz0x8ZEcBAnoPfPXnSTL4boTw+SVurdCMAiE
0K/sTdlInYs6FTaOiWkBKFOb/OSJ//a3EyOlsN7bZ+vax/JMMip5zn5OJSitTd+L8lEKLK4aeIde
PgBMLVaJFX3UKuI1NSbZvbfOWnMPLxzdQ9JiaV941MqpdETg3wacWGNG3nxmKeLxfpMyA+88ZNyg
67quHU2aF0OwQlqh7Q//ADN5Dp7sKTMFDjv4gXAUuzDdXlfSTPVhMBqtG+q1nzdw2M8/Ll8pzSO6
JnX6IDcz3lHg+1XTlJn46/OKGatHtpm3/BvTitiPF9iHYSMjl8odCXQ0WGXcUf+XARzVWrgBIgQo
mMawI3V7As5jTIq1OifvJRGmLqLblT36tkyM5EoRtmn1w2P8MdC4s10HyPyST/MqhFTwjrIfsqHy
sPavZ/XLGN6WSDz/m3J3omzBBshceAiJ82Pw1WyAp+WtUWYMY+fLrWQDu6mAAgeL81NJxMMx53DX
B6D0UP7XmCEgp6uBq29lK1UYoW6O6vAncnrBdvq8o0fVryp8/SThdbjSjA87Nr55aTJjL3CPu/7e
rr8U7IK0xk4AIBY89ZenJAxF7Oe56pv5uBWAp3xo/xVHkYjyztjJc771LIauPwPQ2H53b4UvKlP4
6d/sMCDFLXbZYpNrUFE/O1BdbSNVtcpzsbNB6jUUcwwbcssQSfW0bGmMmp9uR7CTj+LySmNjGeaN
Br9U1zFu5lVevHakV6xEtyvM5awMPSfVld0/OEQ4jh7/3WBzsM17KohMuwdbieTfs9mjCMFGVJi6
0Lkl3iQnuJIq24AlYN6XUdJxRGajAWyNv3UU5uYB0TJWazEY0chUD+AlvJCinU8wisVJXGXLtoKU
QIsqgh+PQNIF9bQPMZfbgPcqmCHkLFasrYKGFlSHHPGX6ENI9BLR1jXgCuTAOj41AcS/6ExUozD7
tMKjPLD7ePz7++FTA74eP/+6/aqdkfWVSPNdcETabiB2Z4DjP18zzA3SgWLJFxcMv0wmFhyHVu1F
zDbCRhAKFfm4F0E//aFM88x4Paw3rll46dGy/SoU1aWNf76uKcBM1/EtiKdgLDYrB2IQkEGUEM2r
eZma7DsDHqjb6NKsHAg8KFxAy4YtJE/yEkMwDoYwHefhnWL+FOiiaxi31AF7Mk6WY9zICmN0M66Z
KskswBJ7zE3B0+JkKIl3mmEWiLboLmUEKhYxi9XqAOpYfT270VlyW4e/3UlJwqUvF0V7oiLx+1E4
zAfLSlret07KGbGIoH/BQILes+Nf5HuTR+URrJK6WpCrquUhbdURODpFnbDOFoocEMiRMcuihY4K
7K1ZsdwHKy+k9NkzRJrDmzxuWm2i/pXd6IjGpbxd1rIutEoIwPd58xl2kNERmXqCl3oyl0kijJd3
ovsVkS70mNae9WqCaJdGa9ALsbaAoamnm5iR0YDYE1e4DYVC8Rp8GAHjiH+EMB0aZuLFJyadcqOU
YojsG0K4DyQtH6pd/IAP4bZHboC9QlW97d3EPbzkGRHewjH+qW2sg+FH5rbz/vbeDGpUBbxnDITJ
bXlFeR6w7ZmMeqf6xdE//1w4eP7eJNQy+cygKt5kZxxMyxsR7+uP1O57xrlyt/tilq912XqXZA95
2bulcRGJ6G74PKvqLx66Of10TF9y9BOVoNbYLJrr/XaGMtwYZpdD/uuTbbeUq8GSlbGhInINMEu4
ko848XWt6PRJZUbR5dc5LkffiUkXzhGiKy9EFicUO2eeN1ArBNfQtx5WEhVfBoxxhCune40lw7V6
g9q6SBtKjKLGmQIr6cWidxgy3zcvMvrKo9oCVsp+2gN4f3IlOKBGVHlglZww3qjvxdbGx6mO+jVt
u8mFwCR10IDjxhC3aL0ceY2+kgq9Hmdz3BP58nbvpIRGL8xlGiDQ2kG+3NMA6sz8zdoL1e7T0CGA
ThejIAAu9dz5X3fG1AgDKO9kzBkh4x73gUJ1VxwBSUGH5Zxn68P3TX3+I9VehW02Wu7e55bQpyTq
FexnfwatnLkGSbUa0SxGSN+SmEL0Eih6fRXm1Vps4vGaHgOe2kl+ZUa+q9t/NjPEsvZrw5HBC318
HNwBD1fK4l2GyhztJD4FfOCPr1ti0YUZFa5/o1St0cG0ycx678TVJPZVd/5+eTRsAACZLje4pBb4
k2EDTyQuQp/n3YWyrAD0Ye1vJpRqpG/4roB/31x4bh7KJEXUgOWhAmkrUDpxkBkb3BUZHy88Tohq
PjU+IhnIV+zNcq5u1ubDQMkCskmgfc0RIXnqZZtnW47pv66kb/PWzP1W4TaYgIUSXstTsIKATXZP
ipqb6u5ftZ7SbU35gZ9AqSpVYC7FhcZjI6EarKRbvsxRw7xhLAKofrHbQBa9QBNvl8bTDBiyKW5A
6AjarhcplPA11m+TPua7f03NIplX5WmTApYYITSoDzHtyUZnVvfmmGmFTe6fY1CLEwGx9GCjJOto
oUnGEjukQQouPZJ4xi1CDF+Gx07YamPEMKQdryk0Zm1XgiwEVVUO6BnPSCkGZThn5gFXLz8wI3vA
SjEniJy09RYIItDwUUnx/M6TemFbP0r/15olYrYP78mPyClzSjSirxtK8g8yH6n38fKSgM/GqIDb
jkFYV02PJ5rVvvUCtBbun6HLM5LLMgWXNfKE2x5Gl9s4KwQlWRLhhHVQbSbPz3BthZyvQsd3E9sX
3KVtX8RwXjNhFSbNFZMWgX6qZS02fVJHAnNfDJo9azgASvzACljElkdTMPh281lM7n2w+qGNrKyn
zsRxFh32r2ZJnzvFF+r/2LzwXROZRj31LuwRzIXxfxjaZQAZWeFl9TsmT79bJCIuPtknRkTMZGK5
AlLK44rG+yOirAw6wi8RHTsgN0esfrJuyLoWGqtV3z39b+r1v4ZcK4vH2e4uwt5t+z+oK2UHWwnz
NYvf5hNo1AlT5Mly4LcTEzYll+KP7B94+VnqTCsQcMMD5v0U0w7+14zOQ3sTYVeGyQnLw7YEoA+u
zir+HixkBrV2nQdo7XeHiCCl1YUyIPztzx8Wem4OE+kGKDAC3cAyxngiEhEZ6hfnMg0iKF+ZHSc2
vtW/ltlZ9QzodCcV26Q8KEAPz+rxR1otonjv7aWqGgbOBfI8ishSkwuwdo8CA6m4vhSwJg6LpDOa
k79Rn+EGNMqiH0XrGSCVHHedxkcAtwUmo5O2J1+tT6D2uF5GoFZhY6mrCDhBg8OnGM6NoNlvnSEe
JVxadsxalGnCXLsKajKfXlaW+2Xv63d8wzf088N3zP45GUoPOX3QKsUzTN4rPcZuKojFKEOh52cs
o6G0AXP2MOpbuVItxMhPGxXydRsLoy+vCZdgOUg64zB7jla96l7sDl1fnTkbv9hz1uue3N07+CZU
r1XRuvFEOFM0MKLvGAjLpzowwBIvYRbDw6e9LG+A54iTR8yFnQKf4d+/TEOR03jMHNE42no9psRU
Acg3CmayAe6HkPzzylmOyrfNL4pQFxDxg4V16SZdHYwSjI8bpc8VANw6C2ndEdyDdTdT0Fo9w7Y+
aVqNEon4pO3LBFCGIm8MeBt1wVGZlhYoXJpJEzUebp47aSRYav0glVtp/DmXwmJ6O7myJQoFvIHJ
1FPuyDDRTclyQ3Pazz0REziMNMCuKz0pCbNLnnTjqU5kZpQZ+QTXGrE4pSSqMZ7imDxUPUBN8guy
XN6giu1dJou6zNcTX6B6aqHD+jYS2dlL9aiBDjO+Kmg39GFOKsHYkJ0mKhDI1wryVNofyGlYaNLp
OwU5gYV79406UIvaC4c1VMWNRstI9rCJsi33wcFnTv2cfXn025PPuWsIav/Jg2fryfsBcy7A4j+m
sQfimgIRlGSuSn/2EQX2ry1ucyig1xAfQKTts95zRIO26htd3mSg/+W9SzMXMwAq7pPM/3fpJgDP
dzeDrpEUoaYFNI5sNk4wD/4ZdBTev4DeSPU1n5bb3kxXv1m8BskHaawM+HxRNG42z4KOAaw4R3Gy
WqyIyw4mVQQvAzG3eeH1012ygT9142H1RvJt2PcKsz04gYigN/k2eKfqmpED4eAgQUHLhsZqzoyI
+PiBdcQMEBHZ8wUcr6ZGkw9qkBdyF4Xq1dbEcflgTzld9SdD4sj+k4yudXYppd1GV/SUOWR/Rxsp
xtsLr15R5gjTZe+hRf4qmX7urEnZ8qwdboKzQxx/hIw40GuCIy4W815j1pppkOno2OFoAq5WxChZ
6dfCXVGI2B9jTLCrcs8rL3FBHsfn/75QVVcKCzyENXz0k98KwK1d/vN/beJMwyIp35o/96rsMtfB
X026rEEgiEToA2mRjnw/uGklRu9rN+LAPtTkDNOX057BUN0sShxtZytXqG+V1DNfgv2cSah6DuUX
Oup+yjIYEon2UL0oO6bwW7T9qYTjr/EBv+IcPnxR+exLxN1mxw1LU1m1D4i4oN0yo3x8d2aLLiYn
NIq6n84uy49jbN/64ApUvsyZCXLpKzQHhcVbuPxVZVSgkPMfXoEFx3rbCgRzWc8yNxD86xDKRVAm
6rDiU2gVtiVy9BeriI9erCzmrstrdyHltpKS2UabEWr8QSqmVGcyWxM0j/ph6sM8RgPpQlnGbfaN
m83E4mgGV5DFTTL7hwS6OpOuAT0JGo6AT/uaG6jMqIs4djPSur7SxZFUUFPSswk/kWVwHFPN8PW5
mLBMwEnIIrrwB9rM60K2s9xRn+IMQZTR1oOhgWpbpJhilBrtRUzpecD5XPeQr1NxL9Mhg+1HkPc8
wcVSPo0rjNQfaXrfM/juYqGIjBy0HhOyFfZw/SjB962ybZrAWo+Shs2iMMuRgo0azVnmr4bAPrUZ
tGVuTIPcRfvcnqgI3TsyqxSVQS200Rg2UO4x73DOHz1+DPo2ZOfzCOwfUIryxA0QpbkepYTXtEbR
vIBNHsLXOa+Lth94OEZjEO4IYzpGc0UzLz+DlOafF1PrNrrrnn8OU8DKFje4juCJXmN9q0etI+4t
H+W1pGgJ895rVX9jU+IdtZqDZxzsKynont6MwO2NruyKZXstATA5b4rJQ/M0Nv1RMvi/hpXZOgNr
4pC1usqbNAEcMYmVsbDYycEUgfgbFPnERu+NVpAXhb3DbyyPUZMClB69Owu5xfT8M6aTNQ7aaNZH
D/nsdz11l2Ad5cYNHkuftsq+w4DbMYiw2VqsgAP6jGPHWGoMOzUc2iueFcduhjVRDs9SlkzMVWdo
4to8AbEMgNzhEpN1l9xcXC9Kx+U+ms8jnGA+Q4XMXMtVUOK4OxEJBG7jxfzM9Bdp1sSeIHMCtiQX
Zm/DYblVrQiYhaA3qvRTFUpl96t/Gpd2qius0kdyXSkNbCl+BU5pksxDqlzNlVGo6QzJUBqo9xBP
/Z6DwSdB76eWVp3hoNkZQhYUiQ4GVGBvItjWWnYk4bpwopjfq0vFcgldF9CmGsVUhqKTMAWX9Jir
q2BpoGXaQiRLqXpYXieUOP5U+OhHK6dOfSa4+j966MyDx3tMYVWV5YLqmPWiVDJUlrTIDB5aOP6Q
I9m9N6C5G3tLEla/6DaqpxZxCoOa9GUCHqseP8bsOM4vVoQxpUAQHT7Ji+48qYQzXaMUF3K7SJLa
8qdlUwfSPF69jFsylcfJT+kSCjmMCmYBYjrq3SjE261/VkccdYIDoyauMxiVswKnGChl4qH2RSeP
QYKKFP9A9ZK6niGr2UnwLpgKW2u843bCTJaQ9xU7yd8DUTrqS/mrPJVpIgyHn91H/vkG7RZt1DMq
V0dqq4RwUBndsAk/ork3Isdme5XhXopC4Wg7cCadw8lJoX+djmVKVqW9XSkLYzPlqcLmMp6c7IE8
Fjwp9u2KeuO9yyeDMd6KzpvFk9Hc6YFB4ZQEkuwtN8lLL/9jwWtbZsbydgmVxQBgIiz69vNFJrVq
60w6Az5NMhHlaDzj4QFF45Y+9VhAhkUfv2YtxhzDWTeAtDhwFdckyW+gsFvvdxNlN6nFTM5VyOHp
h0L8ZMXZijVYzOsHqTsIp38vcBOlMuMckpWrBz2TBGxSBYw7lrRlmsQZFHpBG449g8tkwitrz/Sj
hjctJqBIVExoSTv7zUDjYzNnsZ7pdXbozDJE6YWy9dgCZQchswwMCR5NQer+AHX1iHQoUBpquwpF
mQHuzkoVdEb0wCvfBlusCrDK/CU0iwzQt05xVAm9yiMFd61jpwzNQesLlvmQLVG7pbbPAUIuP8v+
V3wfxB7EwSQLLJiL11FuJys1LPT7AtUXitbkvw69Xx1nHiSGaowTSBaeEIfBp2XL0b4yND8gSJ+p
YhzRRcozm/ylf+assZbs/Slm1F3C00e0tKyg/5Oj+DEnV4JnRsGAQHYADfCBVJu3T4aBC6p31vW/
rgQ5ufOcK/dX4dghv6Buuyb6Wt4vZ6l/7g8RQK+p/X+/yRz3F/2xKTE69BEmEMIKzNHS3s2aKe5e
hdYjUZu92VV/nABC7TzCGxaPp67SG5HZPFY950WXsMMhJ9UNZndp/Sq51LONDyeuLc+IkdkdXSfM
45ZN4pdC8KfE8pc1CmU/MFAAN4AV5Cbr65eqz7VRmaL4yx86HuIODME1HHC7N8C2GXAtGkqASW2n
d8i+ZGOSX5oXYQdyoWiSpfj5z7jz3ZO8IJ8AGOhs1UasFtQU7RXEzCnVwvlsTwVuwy9FpGf7QgzO
e+byXzZguNfl7fF92asdnBVxLFBP2ASQn2XEFOzlqUmwoP9coIOpGRo3IO0L1penmMK9v3vcCnKZ
LmXVY0sKW/dUbzNEnAgx+Brij1yTXwK5KsyklnGPN52IP92ev+AkLwXoT/rI+IG9DUyPsSbrL31U
lDoMf7Lq8t7emJSG28PWxm+9Afoxp7uWZeI9OuZphyNVqQUTJCzw9DQMBrf5G2yUawzCyNnKWmy8
NxxjIlUgdqc5UFshP16P0CqfnUtd7ZMKwLmmhZfchn7Qc96nxET3wFUeQtqf6flKDinwr9ptTpOA
fK+p7Ht6apyfq3E9gKkuZdTHeDXw50jR8YuImfK55+2tu4B7ibDeh+kOkRNU1TvZN5f1Upp81BLi
LsxDxPXwjWipfcHUKhZMyk51ltgBXlGIlptta9z+ZMe8gU4BsOQa/r9LNsWcIm4NrEvv4yYncL+j
yxvTuyBmvAE0bxOaBTOgwJNiOFmFcoFbBFZGmQE/1ZyOGFUvHP6awcuCqPSepNeoClAVqpIVNsAg
XMdc9F1Epj3d/ksY98+aftXTFSlvO2ZspMxQyzfv6DcOhEU2/CzoXWAoJamQeEssfgwJDR46PkqF
iBVtzLXQuob3RalcFZBJQpBHx1DiWzQtQAY9GwdS4hwsD+HUkdDi7sUbAQp+qCjd9nofJ73k1Jxq
5VucJz/QjwkC5JBBjMbXSqmpjgxNVupYn5SXZghE41WbsJulUB+pLtsQxAHH9Jt8fkSxqluK++le
O+lwdVIdsw4Eknqcn5cdut9OPaXi6V5vsEgkAjgj2anzCy6oAhF3AxvbFZfiLuPT1htKCYfljWKW
AZc1iC28N42lRGC4t8P8wNw0+/5EIxdV4LnHNoyFuHKE6Rg+Nztwv0VkTdtSF/MQKIH9yPX0wk1E
XLS0GJEztf/95VLO8E2ugYOu2UZtqYH4+1Wpg5EeXnLbJRjnZrNGpH9XqRGHX95C1WisGeFSfeIN
tsveufNC5qJqJ2j+P1Ns5ESVlBy0gJeiUjlBQ1wMYKEWos6zIlmQzppgOQPoYjmDuZXel1ymwMAA
UHvjLN8KEu8+xGDaul5FJzvWkI0Yk7M94Mgt08baN3FOaptsdjGS/nT4NglLa1JaAWIPEATNciNk
R+PA5HMxvrdcJ9mAnaS8wLmbBFVXhwwmH088nDk7eOHp3SwYrUTKPn3Bs5LeXUK2RQ0pR5zDJwUZ
IGZF7Nc8mPPCfezDIafuBFmNwvbBRI4JpvIA8pYceGRtN/eeSLvqmlGxV17IOAI45pEb9ADSrv+x
fjT6bsEYXYrBMIQv9VPnzFAkttj60foavDD0H4BGoFPyyIP37i93BzCcdKcK3hV5Gd0YXCKAFzBP
/oD1rEK/ckYLyqD201EqnwpbSNmJ9wEb2nKzKMdkNT/MjemiYiSIDVn6bGsU8m7Kk9zKwJzIdZ05
kXYC6NX6Q9bZf1D0BLyAV/XZgCIQReJLM+7rShudmEZy/1Zibu/hPNXjwEXh5DUjgtGTKiW1kepg
iS0kJ0hnIYLAfw7I2fJBSiYhbArGUIvBTiQJZ6vXXYK3azWcyIV1bIbYrW9pGjSRPyCBLPjeVlC6
9iYvlDkb38/VOV3Gs386jmrh5PQtu0hzba0KRpPNk2tAlST92pypYPqvfHpHcSsf7qCyHVsnwM5E
KimFaQ/fpScwnE9NPEXzseUkAAguQpWX8kSuZ68qvoDz4Mnx3U0Qe9fsCV3EeqD4IZRkN64iRzPs
m9Dt3D6iVu5ISnX14R0jl6dqlfs3tTTXUEJw1bZCJ4eHIP1CRG5LO9g1/sZFlOWHsyMLhBHY2BWn
VeKIHRyco4gFCgONfsc2oWINHWi1ML+3VuVJbbciiAaW/QZZ7jIdoYnNgUZwA9xyXkyB4MNQglp/
of/0jKFGDT9rFA7l90UiESV2fWA+yCaK+2fG4spZJ4+ae8LQmLeKl7pZwC7e0z/Su3RE9K+eVh9F
ZtGzl2pTqk0HmZ/hx1lMmiyxwckEcYMb8LfoCGozUVL+KKnR05pkAQo705KsGdW9e5zD+JriT5aM
qjfZvF7vao5B0Vi6PrZN8qPBNj9CV8MXYSCp7+eG5at/EJsnCZ7u2wpiL/AiybULQHT+yGub0KFr
WjG+5JxiNiI2CfWcNVX/EW+Z2oH+SIlbjLTgQ3c9m9JBuuMYh8lEfuMlbtX38c1aE0OMDKB1mmXS
mt6/U7JsSk4P+wNqqsLRw+Qp4mGlyph3GO7sooX7BT/Epxn+W4Bo9MxDtlc/grlFyTPRkTwHV9zw
a1GhHP9PZYR05DnNK+vHPz+FsFvFNEzsJ2+oOW85O9Kcn3ax1aClmpSqtFPCF0G5LKd4XAqNYX3J
pThNGIcEwgEHrS3+hPd/rVenzZHaYEh418KzetCOOQSxPuaZ25C1AiKZk4g+9wIQc8qA9bbRQmkm
FJZqHmN6Dut9qbQbUaVcQnH1fIvBYjVG/PzNxzfM2tp/4pT+4ee+6rPhYN4nA5EmzZK3dDSHYlI+
LCoy+FS72pC5KW1Y9wVpySIxgd17IjBc9oRs6grPOAlCcfr25L8dOa+tpOY99sBtM1t0EZ9c4dJe
rV8fTl2NZbZVECvDZmix/okxo/z74ArCLu/3C4LEhyhS+VGkJcY/nhLxK3Gn1TdrNJuAngGsgrkU
iO72sZ3htju74j6CIhdrz1UwLKsdXgP9ibkn7rs3iCjjcjMQASPJFCBsn9iJ6lbswCEEYjSEI4w1
YwlqQJzxYFPsxDYmCZ+VNgCjzIvPQ3hnoRKEtGwBrGxIZLn9kBKY/ZgSRcaDBVIsXhwrESGw24z1
e7nDyVNfng88Uiy+XlmbEt+o8r2Ecaue2wG3AyAOyjznTl94k0TSvjN+zyrPS+Wc5QG5eidYobVJ
Iykb/4nixyA389Upj/hOSiJAj8vMd13yvgmdN6Qf1CWIRZOYiXMMc/MUJCHJthX0IGi01EFZ0v4d
I5TUeFbu6QA4otDO3RXKUBoG2kQSDxgHvzj4JW2bZWLlSqkzrteFK13HwK2QPPVmQ064j3aWGziC
LMuE+WgVLUKKKmaYbAOJ6EXDpDMf973ripwMjaiCZrXLSKCxUy80qdMAGidNraNrPXuhwrE8VhB+
jZcqpRA+twn5mKON2C0xU6yJB2/rZ71GxLFLOy5d+/vbbZJss7gfpsx8v/RN2RMiGu/SCD5XCs6a
XpV0M9fL/+Md9iuE6iiiEP1cuChW0ULr+y9bgr5P7sHV8PzI9AUhZiOoxTPoZ6kdz6FRMrYKI4JR
elf/p1PvE+Lxk0cVm9mSqyfdJCk8jVn7b9Nnwg+8AiZBTBbAeiWWG1lWESVB1oEEix1odoJNBlUY
Ysv1aD//mH7pOisK5uLmzo3YZc4zw9MDXrZCTJ6vTZuZYQui7Ypcy8aZs+wltJz405Up/GI42DmE
EHzhFapLGNOcJtZgIzBXeAmAdB6tPYEhJlofTwNEfBMzIM90y3S+SFn+X4rACLtkvtsdFAm43Oy6
mWPcSiUQHlRwN0rDW4pwlBlSgtZSA7nq8QMgS1chF0thKYmljGJMngHl7fDILAqnnlTZrIio+kj9
jN/w6HBIhB3hc5SZAnoTny4HKS+i3fmVNAfvmjBlU+TVpe7c1N+aN4tP2QyIww2Ows5cex6HSjbj
sp43gyziKWm0+roHbR694AHNjezYTjlrSTb32IyuodXlLgS+k4nv5f9gpo+mbPzSOG7j9Sm43NB5
AvbgqE9jfy0AsdF86GmURp+a6D9GlT6tpznN6NN06yRuj9WWDIu7d7VS7ocxftvcW3vp1xwEsuP2
zrT0bjbKHtI4Sc5PPqJlXvfNSERhXcDoxy64kMacqfssuQg9Cu1RSOqH0bSznE1h27+J9HMjYqRW
8IY1DqAEMhsigN5/TIkeFGA9wbKK614RmjPFZH6qbH8bsMjXAh1wn5VyCZqc8Xpoj8h28qxkLM/x
6FvCyDsg+rW/WV/zCOKxKl1G5auQkCYo2wVDS6nQEDN+aNnZuBxXjyVlKLPdk+CSmNasQba+bJ8D
QjL2BzjB3cBCcjSUuUzapBWLinNutbOQs566thdMgMXiJ3seQQSjMrqPowsEbsM3s/oSxz8VUQTB
UnpOrgMPrxaw6j01jY5efBMWaf9o8x2KFKsReRtgrtVzM3cg9ug3SbywI//jUvsnf6CvUriU7okt
UcmWfwDPV1o4dxnWDrcrvas1RCVQjNefulvCPk1ZWOrBwBCLQUfBl24bNPGYwb/UiNCDu9xOXcg2
GGam03Ad1VcM9DDobXAsJv33SiSMC5xarkVa+nXxNfR2lsQog8IsMB4cZQj3dzSxdc56ZQyirtPo
Pbiy39x+LdbSociX52iNNJ7mYiWvNExBNfDmw2hMH2+dBgT08JTMuVj004thY6Bc20NVa8AXFMGv
fuKy22ylEkNMUy3ueajTajEWcikMfkVJPtMgsbIi/K4Lj3gMHJ/8cY+YTal6gvUKF/9IkrvCw8ms
7Ukj7SKaz1/sTWpOhrsruUDrNiwMarh2VRRK0hoM8YIlC5BGZWkNB2TnXqCsxiDsEt5ay7jW90eq
lqnKT3xyCASR5Jh7czFoskuSebs9AwRJlT6c9nibcybfcJnBJ70IC3VfquKfKiaMbMLj4DVHd/LC
ui+TiZBx+WUL0aRMC8e8QrMQjTHaLltkEB13VwQQo6S4IYHZ2fdljOssKcr8S+Zqy+9NRPTr9GRl
aVYDCxEivL2jFuX8QDP4Wd4PBW/J1mCK2BmR3t1X4e77/6RESsHddLMu+FgcBCCU51JyGLWxVg3k
StvBJBe8OwFfRtLmAd8A2l593uZFiWorepqit0h6DfpZWWFGEJ/odFRPFAhEpM9aaqg6d06c6LqK
drJERNSj5wCVyo17Qb6rCCDO6e8cB67nFHjAFraOqkm1lx7SMlseb/AT+084MmApJbfGmr4oVrQ/
Qh2sCTJcuWnnxcZeFkrxi+miiJgSSNrkNUXFmKNP3JtAisYGagl6LhmSWyPjArgM8tPchL+p6dIM
lbm7E2909UxrEabMFDxGfrNL3PoltP/01gM1jZ3GHOjLDM7aN741IXUtbr3ItEvv4jekIXk1vYnE
aadfP+qiw8E2Gdg+sWw+cCezxqA52Mi/bWPe00mDVnFkQsONN5ZKU+9mT0YYZ75HLd4Z4q01nAxm
HGdoGnNnSYdP38DBiWIfmn8A41EL/mv/QTrT0hCxogOmDTOhNL6Fs0Hc8KQMvQKFpKgF6OMUDl2L
1hwAj6gsvqPl4OU9SwJQcfWYmUcDn2Rry2tdjwjB4W8hNa246FvLhig0wIVZODeIWyJBPJ4erEKd
zRAXI87ZX+bWl7UTpPQ/h966DMZ62/yqCSM1c+OilELZ7Q8fmQBiK4DxfUM0KmfUHHFJxauIGn2A
XVTy8RVJrQ/7sIaH0sMhTbDY10sRjbSc1JOtTvu7mADCrri88oEDb2ssvh8ydEuNIQT5l1NYGhU1
MCfCEEHemzSu0pUoLuLgBu1+pdorbO3AZ/3YknSoANYbgfAEdMfI6ctZS2jK5g5Qj5FgyWH7IKb8
BX7uofQmVhhtSXiVuNAByugaHkPx3B9SapK/XOcNNBkIelJWkaEKzdRhHRbVmu0eMW5TCm+FzYP6
wtbSTRoDkaP72PotLJfdA14TpIyNRW1FjT0SoHddj9DiWXEF0fpxu2cG6mEGayKeloi0g/2PSdfT
dXO+CV+UnHXRGBZCIfuUhnzrP/waVUWaBawAr0XEJ7A9MAXtvma8IOglwm4mO8HOZpZh0zZavrqu
KPJJB2ZW4Vse3M/cPPJVAvH43zjWgT60kFrqKraktHC5YuRYB4Wh5tk4G1umJ3QkIyGgLc3Iue1O
HAr1NucQ1tcgMffEsDTqizX9kn0IkSz/nxiozXwkBlaWrHWKrP0uYxv3SQTzmMKzWHUYt8QVzX6/
oNHwYy1W1pTJKKuLeIL8AqNFeAr4smYvVoK+KDgOA8F6Ut4JbZxcokk5cSou6O8/n9xHp+1vxB8x
MaBoKLueRYGqgpiWSm5nxzjzJvUQXVskhk48IX3nPuhrM4CrAftBpiyWoyDakpX5/tWwtW8jCZeB
gtZr6I2kBc3j6rtGr9FaWhmVZfCwkeRttZTi9I1D10ndJgrgz0VaR4uBeacVI9uFaz1jWLPyA3sg
dWnk3fsFsuqti3DYIibZcuke1a/m1/jrbD2H6Og+WpkHGJ+5i3LqSP63Sx+Dp39Mk0C6fyO11iWf
YeVqxs3UeUf5mlE1nJjUmtSzmBZGMCyxVw/kXRLswoNYCKjY0DoiqL6BE02O7NEXoLyPDRx1P3Ua
hHbo9JmhMQneIB5bfZl+dxNG+BXLEQ4itoGEh4Ubh3IBL5iPu7Da7MpoTWxv109ddrT7nrbq0LrL
8AQpfjZGzNWqqIFp72Ww6VOg9gjUVdg8oxEvqdCQviQRt7mL3LY+y8RpJ/rxdXizA2ldE9lmKJnX
TyolH5pZagNAmA+H2o3jQW53Tbh5LUFIvrfe/qL3KmX7XwVlGIXIgwH5E8Hkh4sOKQfT4K/tB5L7
aoaqcc1IGi1B3GAWlzB5U9qkHksKpwTOrlyKQ3xmWVm0ioMBENcUg6QtCmhI0fNG3nth8DgQUJn4
ILuhsBHhzLqO3Sk80aL0xQcHW7euMo6y6O4KPDskQDw7r81dg4SBorCEfMt3TEIChx02NYnzamC/
Gt//hMY4rPBOx0XlhgfErCxz6o5JWyBOpjzc6G8RSTFjKbWOGsJoAtnjZl6r6SmeZXkvjkffGEgw
tr5IklPmUpuDae49/wE/C1bnrviKoB9246SMRr2UyHikjIZkoITgCOiLECRCuOiEKnFkK+ZET7N+
XBqcIABNyPcdT1w7mrdJZUD0jiut47RVBW6JsMRKBp9W4KblKl3l3yf7lz+CgqQ6BeuK5+vMjcco
bYwspzEF3wZtcfAI0djl2H1+Fmqiswx6nkHhIe+BGqheEQIy1Hhqeq+PACcRHr5y4EJpir5Hjzvm
n5QpfM1HgCF/s4iAQ0R8j8SJX4b8PJWE7fLWfUfY+2ylcJayYtHbOm/ejaqtUcGMVhtPDEKH7kIm
pQqYbYO4Nws3zn9PZJeiHWBEjL/MZv87abNLxgEk4cnuDQnMSnlojqRvvrXtYlDBNX8tokkCrB1Q
zsDx7uIaMyrXsbgJtHDEYamEYg8tOj1nQpqyqLh/ouucLA5Vw2kgpv85hbHyez8/Ap+iUzCjd1vA
ctobXdg6APUHWUsKPgnl+FXS3XJWHJo0HwFzLnHc71SYcPjwz96mnNARnYbhEn6j/TI54/ValBxI
4xsYF1QwxtOWz2L7otJjoHHsm05tIkdT72BgREuQZCW21n+CVrUu1xIBPLgN3rjVU3NXB3LFO1/p
OFaWR5OvGOZN01ySnRvNBTwdZ2zj8NeuiDUnnPb/4qOkKjK74VVHBFW6abVfHhsqyn+qZcNH5tJ/
DDP73fcpkb7JV/RD473HQGUBaIisp2JZ1xSiFZ7ahQ3Ou2rapWDaRd3giBfMERLuABI6S4N99ew1
qr5JrkeJy2gUa25IPpKX1vvZMAvzPDuvXMwUqM8O7NOagrujYy4vZzLz/aiCWjXDSFfhAHepnQ2N
wTUdfN2ScpWbEjluWwRQ48NyUO1x7DLPoA1jYV/9Mastyqar63RploKDX42EpHhgHgdmT/M9ZqnA
U55aCyHcc+Sdyq1eRT4i8vPMdJu+XuFvO6pYfPrx7GMNC0JM63MAyK7xzuLcqfz4+/1j2+XDiGkO
ClQRzKuFNAzU3znNF+IrntllGJ0HxS+f9N4ZKhA7PLat22aZQD7Rg7Wf3glqiHD+9g0EbKW/dJxp
qbiea14j5Y2tVuBXlVfaCx033/nyYsoUaGlpho0CvCV4jMxOs5NGgyYJUXRjNy9yzUkJ1ECDVdH5
bBSC5myEtf+SiJTI4S3b8YjIaSDY/cQPx+kTXQ900y2yUFw3jJrsaF6q6GAJl56qrsC401vpatqS
PlUFBPZU44/f1os7z/P9WQ6RoAQJSVHLl3C4g3LSL4G3g5XjTQdUUw+vrEDIc5m1wBMwN6m3w0Sv
RqdCgl5vWBZMh4j9S6yIrOUnE2qE2iDpjLJzlxe7b1YcoW16tEC2eq5bnjXqgLd2bpK6nhanOEAS
ihZK7JQAPzPninJTG1c5R7PiRvb9XIm3ENWXm2wF0MbqD5U40kSTz1F3BTIvhvBxDos98ffro2dk
xA61mPRN1rV369FrNi2cYAbpQmcRpyOX61fziiWQ1CaxbBbCOqvIh2S+bIDhr0BQGufQ6dQJBt+m
qYquxegnqXzZHi3CIvEaESlo7DQqOns8nv6VrgaIA50zJ7gsVOIcxaKe0URan+3hY5oaxspz8/6+
98NmSOkI0MJmbomYWzkxmfW95Pxms5CrLS3Vvt2GL4GKKaFauSfwJ+Y7ThtDah6unNMq9HhJ8S3G
QN7rweVPDODFA8JQ4CKawfwIq8K1ZDNZXceZESyZOVU/gaBIbGMIHov/C4tAuV+r6ojA00n1FH2n
2ZClLqasUTeUl0ST3jBn3Q0MyxS1SiHZSSSLIy5OectiICI9GWN8xmKEhgC2eXZd/kT0ve48YL/j
0PydlGWLnkLBWKFKDJ0f2kdV05rNmJawibW2tHE1gzQAslb0JEDw7fs2O/qyUQza/SBHuOUjEyTv
ki0K0hkjJNyOxFr6c7aEn62AjTyVr5qna3I8NcBk8Up32TWh2sPtA4ycp6xGtGe7fPNfxDRP8B+j
esgIiQ4Jq3QghmGOL7IpVwMDLsqOiZlt4JXChbcWQFaw70tB5Qa2y+dhgSv3T/z8gvzmjnc7BXR8
Toz+WcmkKqygQxFtKTnij+LOcAHXIi3xoLttLXilCv/bxZusG9rb8/d/J0tBll0zXFJhRMbWsA9S
XEuwDPTc+vK9nX1bbwmskhoHbwkyEpZzxN9oPst3ehHMoqr8vitEwgKwV17TVM7nQVUdSFIWCXz6
37Wa2oqc5g+OnbW0DAESKRgJKO4mO3OenQ1u6RLxU1w15HLwXDV0ujBzlrE5KEEg/mje8urSKMfi
/plPQkzXo5F4Vn04amyHOD+o0de2i7TjMllxtn+TUcYXB1UPJBT4srkBefxse/tkpEva3wOnLTtT
2JLqG76JYPsJx///QcpL/Rtsk3UyOvQ5DaOEdF+Pa9ch8/WmmTt5PCLNqjJQDciN0XTbhJnbPeGN
YAoUgoM2ymIZRpjMhrtK4Vg3VynHZTWymAa5oUqObC6Ip/es5UiGD4w00SCoInaeqSvJh/03pYl3
CP/tGfQyl60ai2s307aNlL94OiTYu2ASD4AY7Jp7HHuNDLPVNYSVPSUpTPlhKFWYj9KrKtZJ31lU
P6mIavgA7D78hjyFMBbEpFLJj6RfT8yhMW28KE0PfRKjw/wTtb/HV0ZcQ2rTbZLtMmekkLURiKau
6JwsbViz5vEwdakvRN49YjMyC4LoPv/m3tKgXua8gdOL4zG2TRTWAfb29UhAcF2/gcyM9oJjJmyM
pJm5dw4pWnGc8sGnBPpKIDC2Qsmx/CdvtX01qAdfh2ZDhsqxMEPox+N7rCUU06Xu55WR+QjYDjAm
9pK7tjJNMOfBYyVs93sXMx5HGy3jRgl3QWOXMvebEgQiDGbqCNB4AOOhiSg/Wo+FnvnrUNpIFdeA
P4RFU30At6KJnokx157swGt6tFtbP+Wg9/dQuOOl046+MQ7CzMOgnLAjYHxGNBc0klUkW+cIayhw
dX6CP6hqCmpk0wcjlOiM8MGov/YKjEScFZa8oyKyFwnwO3mczjXTJgC9Y8Zs+TV7SpcSvM3E42jv
lpOEcluU5QXYpR9NHJSf19N53TrLaLd7jWo90awZ1u+hLhb+ZNZwwiO9wjWqvg7+h2JEENW4voWe
5PTGXWaXHz0oIkXXvQAJBdXpdM30fkN+/2wB9sEem3gxQYvIQWeRGChcZmdunqGgIW7jOtTWn7lP
0hmlyAEWI1gk7Y7tGL3KwiQUMj9BV8ryXUwRSGWaNPM9hLZ73t+LG4mW9012JrHat2/SUBgOwDez
zXGEOLfzZZltkYFzSBnzxWT6/CXXEy4YSGbndTbf7SA9Cgd32v5TZaMKfp+XnqNrvd6GLOAdnbjw
oWLGf+YGAi9lb5bL7uLKKDEajXc2NSTspolb9VL4dap3dzeXzhybO7uN9Jla1ShfkBZvZ7487V/M
cMg/xVf3Deo63hvoegx40StnR2Qk7/Gvc03wy6OOWgNN3nlGL1vmKeXhDmAyyns4RQ53jeDBberB
Z3re6JQlTdDiYmzEzZawTVw4fsc3vsHVNT+6QQnus6P++puxgX62nkH+QEU7+1IwUcWw9c+laP1u
8s4fs2snVGNueVAPJ0tbgYY3odbkDcaMI8GleE5WPUPFHgagkkUBsJXMYiSr2NxiTBTjdKatSaaj
C69yN796KcGKEYf2ZgE4Lhs6n/DAg4L/0I6EtAru1SGpYn38cMSNmGV06b0ynpol46fYKlqXYN+f
WdjXiBk7XKgHcgeY3uJ5bi5ajQlSrxzbBV2y/unGZTZ9FWOIqHFSgys8TxTgYiFbZhK6WIDBK3WE
+guAEjxgELykfKF6XIPPAiUFWAaTGfIPTsopdbJk8gtSEc3zMmqWmiIt4FM+SI65AoY51Cy6tztC
xZJvKg7078C6Zjnaux22OZEDT+dAyyFO2/0GzpxPcJ9q34mpe14pvTTwJ7zahlAm8AO8k1Gfa+2I
7yS4G4NHMH3IhEc+beofx1ymAzGnpAwt48PJC6Yn27OCahLwuoRJZL3/Dxb48RpvW713SIWcvPZ9
bsRNEH6UyLQYCjFrhpnRB9aLSdEXsqpv3rg2+rkDuj8+ddcn1pqDRIrZEemVonts54C9gSbHInaH
Nd32d5FjcDoOFdNIrsiiSB7NHxx/3lVYwNdan/kApEPzN7OXjW/6UM5rkVrurfva7oQrGBuGoXo5
Mk4Z0VHD8mjg+gmsynwJV+CgyP++5sy9PE6m64yRNHFiG0yzsE0rFK3kaCm/8wjOLZmr7zXhp4oK
Tlvg6QuzxEXEWk0FUH0hol9m4VywClgsObTI4q227pZMUElHUkwHCrJU6WmAn7kU6rdIiXPexeZ5
usCwFumwD3PuwfmeeWMr5K/g+glc33bhdVRKBHMnV7r9eM+8iSE3YnaUw9Wn1HDni1w7yHNHZA3H
c8X4cU5RRFVPaeXfOXLtVgLobBxEZNrBGYm3V7Hl0m+08Klwd1KcWSkxvexVh3CMt0b8J7mpi177
TpK9bFMrBS27Hwq0dZdevvCrox9PdloxxI5HuZ76pPHr4oLWoKVPTEyOygSQ0GgIqjuFAz9Kxg+d
xBYraxEhdD7e5eIAXipvJZoST2dLxhMb19uD10m6k0NuIAA1JNUhn3CZVXrdB8nVTVKLglTplTb1
Wg9v5Bcv8jq7+/MzCG5zkIwbFQGNpqC4wrLJ9dPxEhOdNZHadqWk2g1Q/dtALO/70H5jbT887k2x
ufvwqrw9pmpP5UxaghWvcR+Ay2Z4GmIDvA9uaCek2whAe6NTzO3+D9cjck2hN9ko3uPJA/bpGRfj
MQXV23y9xEsb/1TD/jZOzN6EldDKeIurCH5cTN0KSMnw5Hg7rIYQ+SwnvDYiz5T6Hoo+PZQ3He00
SXZXpYJG5bwqKnysudizEMhbPUTCM5QUIiqxPR3pnFqndtVZFVMSoxTf7bc/OlwgL/2YBPi73QWs
LmzmKkwyaNhJ4MW6JkMsd6YGizVEgbi6I/GANfJwj5jQ+/ffsq+5rNWVSzK7kLlqoCKqOqWvlMMe
tN1kKAV2qHAQ/VXNuslPcJph/Vd8y2e3j8BIldEG79ZK7rDRvkq67JMDsrd+3lNxtNoyUG1OAyeO
SVlTeD4tNvBXo82Yq5bnG7v32i6nnnU/U/uKGC7ggWjcJzZX4PIoJw5JpR/fmfOFp0HMiRBTivgg
jbtNAzBnPpVGj8s/dE1hGYBxMwzQSaG+3bSbkZ6kHYvp4ecDudZpaHAVFhSG5K77E7Ljf4J+/xXJ
K/jE96FxFHnRq3lz5b0qCsRq2UCdiKnW3BXm2IeghubT+ljIvtUy30vVomDpbwh+M2P4qXWYQMEj
kIOwtdmoWjwI9C8qDf0GuD+kjk5NSwkSYYsqHyaWRS3SkpC9r89pGP5HVzmEEpfl6ofMTnqDe8zx
G5eJQ4P5/H0QPDWEcr+Tp0UfMGTknisKGWa1gCoC2kX4NInrFSY74boxFHRDCiG+FyMAg+aVQK6V
3ZddLNOyJKne82SqSigun52ZSvdnvrRr38SeY5mCynGoQgdJqmunSY88JiYfPbGE/uGzEwTiOEH8
mxvMkysnUUkKw+u+0QEYFAwbLEiTKY/yaw8Tomunlv1TmGi/O6Cg7fL/tKmEqg9RERlZH2QzrOu+
roWK9lj/v3pUfoKu2DbAuGLgbHOAKIZkbXQ0dvrpl9cYsW3mxC4DzswsN4xbiUkj17XG9WojExju
qdF9oya0r0NyV2Vb3BwOAGcnJxopu17r2SdAOGyGaLFYe2zkzKCf63ZOc10DVfP8kY21gxtV04dd
VXJqlR7zGX17izT5YasPhpqr7RzN78eUrG6V8t5mP37IDwYF4uBS6BMRzsuOeMYLGYLPK5mfRAmq
D28oK9+qkBvByuLir6WCl+kfYq1OX+oj9vtWkG1DeqxbsXg+h9NoO9lNbTVlW13NBpAhJekytSJR
3nEtEEsglQYzPZtBdrGM/L1reXXBmqpa4IGlY0H/MMrbaBiXkOuaGL2imE9L1ClJabqwYxff9gsR
Upy9SMLuyaIIG6/ZCo+ZadQTU+sDUNEHT5uH5SSNd/+L/VsNufYcB0EVGdD9jo7bKvWSW0GVITrC
hBclE39kSiYmjnfjDYfXVmY29ac5QMuHVnVy9zGfOclNZXUd8pteB5MjTOQ3dZozxbagpc2YwEo2
zm1xcVBu58w8eDnhm6FTA6PpsVjm+Uf3c5iN/s8A/Mkk+TKY+egaWYGKtgS2aM91eUjujQQs3nGy
yKaVSWIwtJC+exWpaybEfmGoB0cReZlh2+8JlEW2iTa0M4uzuZ8DSOVMfPUapbb08y6POszPTBok
7T3/qlkj/Zy629Pdn8T0MLTGACbCmxzsBslzUEQDopglQ2CaLwBEmzkhnlokJAndcazBAKvhHjnW
jJ+6Wcx1g4JkCZikFYnTNI2/lrD3/y/WbovWjvgt+HkMYtKYe1mOixB12Zlh2F5KQLBQxo0StU2A
O1vioQjuZ/DR+75dYOTrtICMfLt1BNbXQRo/Zdyhk6HBEmpMX2jRDk7eYhOUWllaEMkVlgZcCoug
tnBKg8gwo/1CxnIh9uBeFkQHU14AfE2G3Yw41NdDcjEailIBbwh+IpzWxrLsHZ55fKE5RVUPejxX
IW0Yi1ATOdVSZMi7abrk5eRQabZAERnnrW5Gf4NTBqSZWd3w7R/up3kPtJ6f+uYv4RUgjP91GWc2
NN9Z4mQ89z6zw9rSnjl1SNLHxK01o5WS95jhIc283KvdN4c1/evzzLPJ1h+iSxKh1TNkhLrx+AsZ
O0iJbX8J6nzZfX+XgH3XLGqUHCtyZHwfUCjHiAxH2ZHbtpS+RKhlhE+HVQQkTdw2kbY/1nxrYQ15
cs0PsVqZZDmrT3djUdfjRX7ZmPBr+Or56ap7H1nV5iHe0qIsjujVn/xEh03NfBKr6tBnpLJDCXFv
/KC9nuN6AH/KR70Ok8ZWp0VH/3d683ZjU8zkpyh7jZn/vvLpGJDtJ/dxakVg2fyvAx+RqnQK3ahz
GHTyP2bTR1Jh3/uilINwWvapoLouBdqzGt4C0meLWJvJ3NZ6H+JM9ffOIpVZGNeQZoM/lUfRs2dN
kfjRTJxtgWsslZks9Qo9gvgRiusgIiwMsjN1q3ehApr5ANxK4Y0Q+5Ez5KBXrV6yObOrimyQdno8
Z4NwCF4jIxZx2kfprRGC1h4iUq0mVuVrJGLZN/ZNfrGc+BKp3lWsm8mEDCeA4Nhsa+6HNFylJoi7
TrahbHl4OOTB44ygDEHurph4aAzlSTOH7MvbDUGqccDrmLhx4IBxAGFX3CkuBcIZkf9RBRLAirEL
yfks/TLnX3mVwqTeP05vm9Qa2Pw0HRlXXg9Ldw6GPPcKUuC79Sv94wiQVNCkxz4Nzda8F8IhRyFY
dUcpZH+HUaq0z5sbWmBIs+EuSXiV5PHEb99vusvm1lN5Mf8yQkcTtU14Uv2LTR8cLon3JE4BowF5
XB8yWQmGG433Sdq78ixGH1qSp3xa1tvLHTsSyxrD7ewcWZyMuZ+m+mjHFHk9L9aniaY3gXGpBUyV
D3CYwByUjwG0ueMqflkHuLJrAeW0EIgF9HDWHgSe2a0Pc3O1l+ap6GN+RsZLSz2mYvHmWB62Oq3u
ZI0IZcpQ19Oav7uB6P4tHQ1RdVWGmAJRubebZmAJ5CZQGsW7nDCSc0aNkleRj6a4FmJGAlaFmyjR
RLZmTun/FqbTi0R4kB8C0KMxTSi7fjpD+4xS53x8cgCUkMYywCaBNJO8UAF91KURXKO1WXdEJIbS
UMy33KvFdGrSrMw11Qg9lbUtAbxb/gsntunc0r76V2ZG1P9Wh1pXmnElLW84md34XpLTeZ8LQFvn
AjB2jwaUbGR/p6B/0/qpbcbM4yzaLavRf1UztUjbBo9GScTptL1rP6hpEJsP4NQpw1OLgOYbgofe
fSrbQ0Oe4VIFWhmfNbJtdYYc8Pbf4rUe7+0c12izQ1MAkcJgA3UqY0KsRr+doajvRsqjDwyP1Wnv
ksfM56CNmY7gd7lB6iOrfIm6adyojm+rnGCCQZeUbj3pOSy63ZtVw86qyTQLQjnLwqhdOLY7i7BE
A5kfj/4vLMAQPN8zObks6+t1M1KQE3biDCOE7q4ukHLBTnb6EnbqvCgdzLqcPLyeXazsaL3wnzIt
o7kO/Kh7JvsPWcJ5QmI79zjRs1NbPr3Tpgelr3pEb0NVpcqN4z1AP+Yg7yvQQj3gtPVIxQj9eGt0
6jMuhODfjIWQJgsk01vYH7j+GzfZWEoHft7V6sbjGxcSCK8jM4GVd6+DGX22WsqWlxw6DenMflMM
txIMKhvckwmLxF7x4SQgTaj+pyZZCp4vuBrttqLiI6WmGFK+Jw3uImxhJWDT48jCnHMgiQy5AQpv
WsURv3j+UFnEbC0XGeEkff/0ZfeK04h+GP4hhHwgY5ATbjvEWgxglrNSeKGwLmgJVeABxNnj66Hf
vrCO5p4n1XR0VHbXPwaU3IxyakdkeVNqx7gWRBlxCbodn1v//0KhsFmVyPOzbkmNVQWkvJihakvd
DJbqEnsF0zXQxkilAdB5TAD0g8LimBzzgathWjw9AKY+AWElvK4/JOEzDavzImxnz2FolmXtW7Gu
drqyWDPQR1peocZq6QKtCAECPciDehtp49xWI56Di2FBVZxHr9geVZPeruTkgWb5X2iNknuYSGep
gm/syw+FzsJBx3Mah6XKvJ6Ogxvd+cn3e7JlFVJHY8a97rg+092NnMN+j18zJ25FxyJRxoOPqmmS
J/PpWPT3NZT6TJMcX9X4vjjX6oUs+aEc1spnCgeBBfWbRT5lDFCDkBtgQlC94CG7K4uIFWQ6CUyN
qgEGU996+PE+5q1YfCBjOtA2YOfltY0/R0r5IMieTWE3cuk5t6xMgeg29ArtN0zpZ0hM5Larr16c
cSAsZLAsi6b+dNaCJ/eMXRB3++pgjEK4LSALdHKZMiVSfJV3GzXDWlv78eIymnSvnfWkNnnn7S/S
XqC5W1rPB6BzIKwLkQ+efx5GepY6Aobg16CTReCkxZ5W+LN5dg09vlZF/cs4Ua+BIWLXxyB/hqlO
ZLymHWOIwvPeiqZ9YFtv9v3w2EatRTiA0Az6y3gnnCIiro+NEYxtkqQw3NzPXyFvs4wXReAXsqr/
UfVHuMgD90rwCDZf7eSgEnOyMlCoSnLXxVSLXb+FOtU2qk9juz53a7gryKAb31kUczCALVsziE2+
rb2wxbS1Oa38n2GJoNkXAIBVsHz+c4zzyELtpbCYwb0zWEQNHRO+aD6nHI3bPU8ISh6KxZ+FCzOi
u17c3kST0nKQTpco2801tKWW7V05iYyXlyN2ZBXj0tz19OXci+4kllxmE0etx4ZwSU2CCzr9av/k
DjBtPlHynw7thgRo3VZ0stMx4D3Y9mS7y9WX3dV7CYmT8dDIJ+T8fHAAreV3URP4shgQ/72DizmW
t3Hq9As1p2hDP89f1H1gcwk6b8/D5HKSIx9kf9R5LyyGDnHHL6X+stzeUEbQGS5gogswrtFM6oL2
K9sqkWY2m6j6JKSkcazR+66JS3UDVlf26pFpXcy24iJSmEOkqn9nUhhd7ZTFr7KuxGZzqNxP39RP
blt5KQINVII2eNIHZZpjRyoTtL2Z82O+a4sXRWzyF/ilEPN2rLEj4WiNzZv6yWSlWhfbv6ztdrgf
OwS0LTvNpq0yeLAZ/xEMoJpAoMMuTrB14NrtNb1BY2Qi0JG26/u0ZNO2Z2lPLLkZCBzhzWc0sZuO
6JI21nOCZo5whebGQsR/CQGpe2CciWMV59t1D6QmAaaE5RjONd3ivHqa+n0yrHB1ItgeD4gLfl/v
4IoV2pZ/IwXc+k2yZwtGR1eXDyEswt/E2ttP405zbq00LqvAtpOutS3wRwYYlcxEbHW4Ku1qCqC+
nWr3EftDLb3lRnrPONQmsKDFzj632NLMUBN/RjOgiez04Bhldd3BS16drLbXZkOhrryxeKOHWxVq
3XADS5G6R1RESYVMi2r/P00FkeFx2d+5SVBnifxNtJptOfScPlbnnrduhYBs/BCKTxSKibfwhsjB
K66YdNj5x9W5lESqjEs7ZFextQWB5Y4xXHtivj3P11ze9TfxHVKKoc8bvCQ9h7ZHnLg62rRmAgQL
ToSY/J5pywe9wRZznUupKkdaZmwif9Z/oM9SqujCnHRiwVVzDM06WaJW6ENEyvZHfTJxX+6NYpUc
XWAtgNL9TZZKF4LNAB8n5tLLN0/raU0ZowzmJ4JL6XNlfEPgwwmihh52suKSU5iT9+NV/BFbx9ME
69I6oIHzJYWah32YX/GrNJRfevkAWy8v/mrh58d6p8hjj6B34Yr/MvqazEXDdnSGz6kX1Ql/xJ9l
UcCliWE96CkjTrIXepH1FVyjkJrtrdSYVTENE4KtAm+kpZ7eXGgdUBHVNe3/az79MKs8QaL/iUrh
RlWNR2Qi8NSqP5pXs1lzW8Won7FMTZddkCQfeXJBqbnV7bvIwQucgFsnW+Mgx9/9RnAUEPEvFz4z
xPo+e/ah6U+Bj3lPAPn0sgkS+4DEB+nqa5qnh1eUcKTboh0UHP79OrzKjtSvP8/iGh8MoqdNWe2G
uXkeIeDyjoJ0sIHao80/VKnddQs1aA8T1zjOenQYlId4ImvCc5MHuEGloS5NU8E75dK51Y9id6CA
0E4cE8igiLSg6xmttv1qXBJTFn7kZPzpSAW/Jb7ruDDRFc7+REfALUnJ+SNPpYSAQrIvhmeq+rgv
jVRr7+LqKK8wuiDFXy49C61P9TW0x9POIvLnldawzYu//JdjDpo2q6M2H9ON4C/3llLgKQJShwJA
GDEd/r6tJ1PoJWJWt8RrmGDFEt1YDeGtwEzr/uyoM4T7tp4YfNSa3ni2pHH1ViSJrDB9lzyCQ3il
fkunhAl5BTkVgZ1iPDsNUXHM5PSXSu54/gDk0bpZfbVAEUsssSvAMyVC///nfa2eUbsGhn7QeCwS
Vqsk5LBmylCTywFWqf2S6jiNSbJgyH3mYzj8kgDCo4R3+mKHYhw3lIRgGLjB7xZD6C6P1SOQgodw
QV0yElgADdbz8r4AA2xxqNMbJ3iZkkm9C19T3VVixHf/cVdfC5fF/QbnBr/bcbIAWbV+Hfd/ezPK
zIv7hcX1KAL6zMnw8SpeE5M+MdcvAC1bN0PA6S3TrHtoesOH0wymTc5i18gaZRqEcpQqM359GEyD
t0xb0KZqaDBPrEcT70iEjDqNnZCfoWuMNZyOkkECMSoKjbt5fkEoVUOKHmevYDffWUr03y9tvcBw
5W30EUH+h6oNinDeHN0aQBzTbnVZOVO12GW2SMPNkgoy60PLQUU7U/YstXfs/jZUaizIe4Vf+fJZ
ij2bo3eoD1iElxWP26RIJjoYZPONAWp6vZ3/S91LpPvUS1iWoL8Ybg5PFvyzs2HpymA6ctq/k6MV
8Esog6MWHQ57DR3QLGUb0PkJGbujqw2BCW75+WNrjBOACCxvp9uGHxTZfKtJrvJi8juhQwXjBXHT
Ujh3E28NeglUwcANjnID5NIJ7TOc68eRbzn3G6MCuOAYTBmfrLxH69dnRo1gEIH5u8PLRCB84vbw
gRzKsajMt/13+gW/xBOZ7gzu6bFpy/kBapAbq+piaBSajR4IzruPUtQPHZQYY6xDyvRV0gL+sFWz
bJwTjrtm6f6sV2PLyKBD9oqVr5bOrJH/5PHojv1XK/tj1vpWErBnnmb/NkI7lmp3mXrUS8i1oZrx
dRnuWZWNyB7pCMNqkg3pV1v2xjT5z4EcCc/oczTAuSxXsidi1w9CYJO+HaAYXyYBO6HxaZbqMVbu
qlVwg/EvNhzXiWIz086NgjSQTCHpkBW6eoriFiIwng/oQ1DGx8dOfJNlGF1fh+XCNly4Vj9B9PGw
QZyjxbQK6XHZmRJutumuz4teXAlOleGxABQD2Izz9N7gVSObbgdptvMXQtQZIMhMLLvdLcldlCWI
rgBTLNdTAnBV3QyMWfml9TlyPK5LKTPmkInR4O88Ns4fleZQAiP0w4biGYjp4rcUPzYTQaRZWw97
0Ml2sHnfiF3LAumrmvxPM8axa/XI47DiazVRmFWMJNu9CSuAII6Y729yU5rZl21VDhNl+jKH1vBx
7I3xCo55GzacXhNY/kyToRyonCGBQVrCZXLw3g9QpgpPtzHJhrkaHO6d0rbJt0ge2/kfqpRhFzi4
8CPSlhJqw+Fyx7kZ+5Yp7NZtVFrmd4z0YIHw3OI1yCmhNhl0j3fMkFThNs7p+kTd+MLJ1zp+Wu0e
gzn97+5K9AHFlwVPJKsDSIfq/cGf1t6y2Lg7+BDd8D83/AufpIFTih0kDRZ43PL0JRCSJHi2UVIc
hFtJ5BVKhTmiBcF5e44lZJkzSSDdDvh+uhL/lEfOyrVq/xJDuKrnG6zy8NEEG9SeyLjCfAkIw/c7
hhYtT+xmeJQ2Mp57iLnRyitFHiOglC+sb2IWgYg1ow0U2lZw63tpV8ajqifMJKmriNR6Q0vz950Z
Osurq5/KvRT5SoLIseQRSfhudcnLu/NwQ69UsTYeuTkPvUH9Kyl/Bhmei1PxvmF57a5K/ZqudID8
tDBwZjjAzmT30+xw8SxO9aAk5R9h6qNxwqm5chkP7UaGDgffzH3V2c9PgAJdTGjXg1lj032L12gq
2PDrpMntdKYnVByZjEjENeEa4PIknviycAV5Y68MACKTC2ruUL7w2uNCfrhVCOKrrTIaE5FzmDuI
Aah1XBwMwEEfvNpE0VJLQUHkD469+hMIWeoQAuna5ydpJn84EjUdOlRdmK/Gu/tFIS+0nCfanwtz
zhgq7YumA5kKsB4S9Dfr9lM4MCq2iL3JC8bYHC8isCoh3Rd2g5DMJPEr7bW7R7EU/R955Bkood+T
1bY7VBPqSqCJHRNvq8UKWeWMk6jIGqCgHd0MHNqIEm7ZJLHvtU01HFIXTdTDtej+ouUaozVj0ci1
zLT7pkm9l/n3lxzY2y7RVk3yHGzjZzZ7XJkpCGAyu6OQA4w9RUfEb8UkwEs5FccGxajhWmMvhGhj
rqgyQzm0Zp4n+icrWwBSN86WKi44aqaQ1OHOjzWcn9iyg9lyKUkwU0RjDTLRT5ErHu8q4KoP1+Pv
/7kZ8zvK7AjOHQWY7BYbHNL58RghWz6idMiMoXQpC8ewSSTlrH9E05h/+5c275ZhFcW+YH74vsDc
9uiTj4HF7gVa9iuYddDz4A+KBPhgPUUlyGNe1Wx4WlLKKFK0jfIwa4pISSz8XWaZhQIvJ8UV4jOg
vCVYmi/iPI4y+i05A2aJyeYhpJFww29tXdGDtm2gvLxRdSh038JaWmKotnpmkjsAkQ/UnMZmEPiF
a2vB1XUl9mYrl/EkMdNbU4b8t/Cqh9AnOA8IYCxnskglK7EMvdEb0IQYzX6YBwIjbuH9QDI6V0hw
rYl0AAWnLu0sqyHxKhDRtOVXZ7wrA+q/rPOg0EK6fMP+cjkPO8Rri3m88YEEYVcIsGW85NFuoKA2
jFqa5CSiQDc9RtWeGbtSkqipwEDH1hzAht9TlnGEfkZ1ZlvZDXwrR2hCBcE+jV+b0YRiUIGKYMLD
7TVOqJPfDTmPYZ6OIF/gE1Hl8ojfMoOvqqQ85tgwU6Thv57gwX/ei23TxLa8GJWg8pMeShYFB4jk
0XWPQ7yAfctkCBRPEPKN0GnkEJ3WTKUap1OXQgolAcvWyQok2Nsp3EN7dF9JXa+n5Ok09zNAZVcr
ZkCq+WT3HZ4xaUgabqHpRbJ/h/m/Kl+FHgrM9uSMWNQGWXJqdn7f89mrH/TX/srHFlbdv6KocCA0
MXvZAOO1xhhOPt41gMpSqNYFf3pkygLJJbcbxSh5Or7aQ8ML0h+iJocMQ9piUnHVIprlg+nqujBK
ZYr41RQPhshvwpH4GkcKmfiSkeEIYgzBkuwghcluicZ6k5XezHJEmBTHeqwYTEGsc4gaNkEt6LQz
iKFqjReoiuBeFHmvLwW11Sd5v4mdGRJeVHzDXZ7W1xaRDXssEzueUfVYS65C/nvTEAI2k11kCS/a
iZG58Vo5yVvvTCPH0RnfejV4tEb0srOntneOOvhUI5yqpSkbVaoKB4isoVhO9nrhGhPutnot1TUW
lp7n9yBdSLQbr+xaksDGfoMYiRANHx3N/jgGkdWjIo1YadMX9oYWxyoHCgFCMFoOkufu95LqYMxQ
zGNS7C9Y0CYBQc4V/dVt4Z5dbdHHW1rBwe6MwDWJnfMPDdg2Dg7FqXGCNk3w56zxvmRD4Dt4beDD
JvGNn3GrSWnYp7U8VXrHhZikMD6FbffOfZMXp5qUCy0yCHXLWPVKscU452v1z6/UhINZT5D2JATJ
j1FtSF9ZAD7Am+naaRRc5esnKwkxXh5iTsZcvn6aS07rQaTiHxrvwM1S9ocxorBIVUSOafVzjAkD
3pmR4HPEcowYiIzw8/0d0Be7YbmpI2wojpc1zTRH+opm80NH7L8w6laU5dAo9cyb1bo3aeuuAnHZ
y1pdFpvvIG62yneHSUuTmQjlyXxXHvf5K/+qYSlqRvt43iNWh307UQadzTGMqAkLvNvOzqqVjcST
+4pu/35ZZBHNwU94ZphGicnhxQXitr0daNXGI72hdBi1WUKcr6Jkk9tAIPGnPc1NSUNQwbDe/kLp
mUJGGkLPFdGDCn0otXjsd9ffDPdJOq+VoVi47iPnzPT8XQolkP4tcnQqELRNgbnM4ctzd820L1jT
W9LgOSgAJL7029KAd2B02k88uo/Bx8yAEs4FEhJ+AVNJg/T7biM6ipevqHBsHnwssd6RhX+Iv+ld
fjj0X8na1UZ3Rlj0sOGEH03dBwITBpjcHS9sEpGEYtXcipaSdHgc7VV76T8YRcDyWzUrP+Tg2OzT
NTZZfrihYoegh1lcumTQ93HKPvbbaQpJCs3Ymu3nL7PQA3FeqLXbTNPTOPSxruwdQWgY3i7i9+ha
B1+7ozFdd1F0u4INjK2abjXTbksf8Jus8lXmrnZ51nFVRJcyE9QdZj/dC4wO3XuZdKpiyHLWjHKf
RDlh1gbYvxpJjjAHmbKR+JOMEt7lx0VVAsNqxSbbNCkrbgk8GIemPNuMa1XawVP4s0z4wZ/eiHBN
np6VBTCMKo+XySUnhqn4C4+asBVWp5jc7l/p/uto00ZphFM0EzlDyFAwpssNz03kn7y8jg/2d8ap
3wfLgMW5XnO63UiEQA5MJY+kd45yaLRBmtLhz0Jr8UqmTZX1IWEagDOQ4TiLzuL3BA5Z7pVaoQSr
DpT0YgWudPpnozAIEO+0IB/B46+zD6OsRI519T32mVhnnVerJArcFw/nWJ/+pP28uxlqsA1YuJwR
fY4fuN0bpx83C1flO5hmIkqqWx2FlCeu8FrD0Di1B6rQgWkPSKWJyX52dUaU8BSn1wjn995MGRkg
qLn9+ZibYk7//Kg7hj0/TXmdd7/5RCEe8oYAH6eDY56XQq/0/A0OlpCIvpA6oeqsuobNe1+/yR+N
ktz+wx6oHfe1k3aG1V1EtomQAnQY2U9RVAF8Q1y4LA6HSvpS5YbZo+8fJvJkWM1UImuC/kItA3SF
xlXSNxYxwpFzYrBjHHVHAPsWLpjro4CyLmL6EcZnWA6NR8l7xVZDt3IC9xciKuSRGx16fcOyNwk2
bsWUpQocF8DuZ315CJL4/NqGXXELMZN41zNHbcchyXqw1vkP1r/yPIKSb6ZcRpwrGPMowUyaMQAR
kmwqtKf330jctjOEOyrVD4TALY7hv5gUZFn4dGGL/CO5NodMoMATKC9NMte067tQI7ysVy5CgSkZ
rJ50iaTX5s5CnIIZvCDqibZ8VK8CfoLTC1aZn7E6KgqRAcQaxfHQjxeiB0TE9Jq2KIC0mXoT9wKr
sjlVFzP8YqkBBTRJyalB5mcVamkrX7DDE3/iMkUpiRYahL+YF4j0+S93CW3KmVxF9NRu4iB/mTE7
OczddzM5TycMeQX200a/afCUZOezRJ+qGIrXf423mF6usqW/R4RJzhPvowXgHHtHYHHr11cPKnNw
pMpm6sjVn618+TvgdIiPuXj+iCTWnygaXlsC1NiCyuzGTbvzVhMvbQjxdYGWQjeIfKgyezNFJLRb
qmXBYBLGF3G2sQnhEuRlJRUUjOJRJitkD1AP9yjvFGkwEjz+DQCvEdaUdBhffultcxW8MjBJSy8j
m3MdiJhgcqYgDFbYXmKLTzKQmIpqHSKGjBwYcqmrmPC6NWMqCKOfergBGHvPXEolBrVl2nALjppN
UzwrJzfrHjHv0+IRN11BblGEaNrUBNuAFeswerlIowY7S5i7gqRDmc1t192gwps7z/ZkcRJgg0n3
mt7xkgGmimAzgHxibgXwqOPx0QPXgrevYY5RcoJK4LuAUQBN/FEhs+sxF8Q2LNg8RdV/QQB0NpZP
VrHxxWx+p8EEspP4N38xlvgkIfH3cS9ZtzXe4uaqlJsaLIVMosThcXouCMbddAPBnQ2KlLwAjzDZ
LUOhIP0TM6a1td2AXQ2SUt/+ie2ncqJ/yyXWskADZD+Is6rsqTCXbxhtdj2ecAyqz+/+g60TI68Q
cmBJgtE5RutF6ivbcfRxPXpXb2/iv/j89PtQaCzTu9V6HN10CgSzxoI7sh0M5eyzSeRgRlgByUg3
tAPDX15dv6EB8KRRNUmA976gbFIKDems0sqI+xqfnD+jc1hSfdMXBP7CJCEyMSAtDaoEuRUFCwqE
KtW7vnw8rE58+rWRGOdWDW8/jU3BT+VR6LtdDC4X6pePjBpV9fWGT0ygb/5XRS1f7L+gjBhHNsHU
HXAEzt5v/CY0dpedckYJRKXkyp+hnun1cGVwVGsUU4nYwgMMcOpG8BqSA7ww4BxYmCiU4BH8PYab
3YtWPaunAhGRYE+S9zydkySE/DmVhUw1cP9QBkpJjNnnaJd8pWbxUuEYcxNgYn+Tzd+B4n2bnbxE
hZC6uydV1Ple2XOWNi7TbE4pgKoMFk/bUzxpOippmVudDbgXT0la2hko6SGELRnRLamGNbR8PJtS
3uGnf/wFmaRrIRWH9Jrq+YCFOorWc+vBs1iPKrCLvGGEPTopbsIj3xSQrgy8OGiwvMG4+v0KoDlD
knrcUODxuKi6hlyHKgzYtiZ6+fdP2Y98fldHL3f7UISa2EQ78EUOj7klcuOAQZ8humNH+r2D+FPV
nNCNZ8+Yw3SQXTq/yNK1D8rq8KdpxAsRmt90LBo1uJXEMKHPXMVgSWW4KJhcCg/L+FHY1UcE844M
QnoxxsoBAJgO4HSLYONYKrMfCy0eq1P/NLuOIPJ8CqyMYjeHX9OF4fF1owuQm3NyPFv/KZeFz+MO
HivYjnjTONPCjvWLiuJJIEjDFZA5FGpNOR2c9H/28+C/Q6V9KRxmPPr/PK8qKfQr3903UpjAy7v+
mFQfq0RECWdpOI3SwD4qs1JXU7XIBh+1D6yfw1DxWziqoTMq2lVqpGtN5061fvUDwRnrVsuyhRt5
meJfzxV2p57NVm81+vsCtZOhdS1NO02BO5ZwuVq1atiNSWGkhwXk/zlrZ5JmJOV5P3eCB2cb7Tdq
wEtmwF+K3ySO4TL+zz8NT/Oqg0HDFexANCLgF83EvV4+5HgLHttu9I9Wmp4Yl7g4dfcZmMIS5h5z
VzSyqteUegpYKLq9TLlqlLmptY7V8aIbVasaGPbkBVwxd7P6JwcsbmHv3MV3CJrBjG3t2QHn9dE3
qON597F/PZV1MwHnzRxXaym4Y5lgK7Exii3CAQeoc63nnHKv4EuEVS7NINEzWDbpE5a9bkdZSqVV
y+asrTGd1GHB84u6V+micLpaWVpto+5VKReSk0abnhIDPMHaRbPmVt/Ah4Z1cYmGun2V/tQqPS0Y
H458zh4BW0y13PM6W8biVPCr81HqOKYNTFFVOdvRKbXoKRdqzkZzlklF7w0LrdbSI/HxET+xYtYT
Tk+lMmiXSDREi4EKrGeBlq4h0sn1ELOhFfyZW/rUWBbi5lSEuK8jGjpKyDHtNJ9AMrAnh5OXCM2J
W6H8tvlSd16muFhrWgMGl2C+MAbrAyI6sFRN+ApILEbWWvMr1qzjKZhx+OYkjs6LhurpbEWDmnN9
Gqdxro/kBDvJlELkjzosElZcbYDKNDyJvwC1UqTLuU/DOidU4Olpcrkj27MrhpqeisAjPGnQWYAY
9CP6F4EnK37FTIFEVrdGc2bSPFflozjy9mxe6C6MMoLKd0WyxBoqlg2pGBnSFmAjkQJSJHzQaSEZ
JRbIKw1a1ARAfCDNUs6nQtft3ZjeaXB6/k2y4eUPEebl3XfvZBAQGldAJk6MNzSQ+R/MfqjusNTD
7x29eDE3ZtPQHG8lraFir4kwsZtJlLeQ9dMefyNWMZLZqyPpqN6bcC6aNj48HPFMw9iSiI5wR/jA
FZO07mtZbyVWnr0GwT2JdYxJngPlUWmWTH2gxXaYtBa3aj0x3nnDutzc98UPyHvOoqsr6PglXpqG
3V5W2R27tjWqnvZnfirD1qJLggVtdJuQzA1W4MB1Hg4nYbtLeVFqYuaYSrxg8jbCM5ASicWGFL6b
+GiM2xu/E7Qro1/OT0fnKHsfGhUdRcjrfbXipvlt0hCZeWx2aw9B/RufVokji+xla5MgSxXJgg4h
jXl1vBkZxgiQgchKVLwLoUcunNGbGtaIHAdmH7aveMRqpjqi7wmtKQ1hS8Bjq8KIlRFUexMUAwNf
28p9kOK0f40lWWOpy6T6F/GGCYQ4aExJxN4sIrWyKASM+yO736p0kCOcZfu81O7zIOqILTLNPxiw
15/oNq1VjOFEc+oj17OKztsjEVRnEhbdlqWwMu3qLrVXCWS37WKriQx7nV1jMHkClMqHa4sT5ccs
BamSoluPp9quMpBFQKexxCvizKDuJMEZG101rVwRCEaiRsxzZDC7QIS7FL5PdJX+Yi2AL947/NOX
2M73S6Hw3pYL110TmLZ0CLOXrkzAZPMVp4jog4LzTYecaiNNy4aQ1z8SPYjnITXZ6vQ2CN1Vlrmp
fsMOQtcPmBKy8SQNdEJcogFT17B23xY31/fSUCtJ0cIjF7sfi1obT4uoLqYg0d2nGdjMQlr5eNSv
+iXpa4edWt+axp742QTuE+3/aujThTNA+HHyogsUvubXHNgspHfogix91VDTLZsmPq4DjmSW1Dw6
5uVGAXNyXHZQvW8eoXsDVS2twW8Co9cNO03DPcjKHj6Rf4vjd/Lo9e5QH5Gwffmf6BvM/jKi3HOi
nNaOnuaR1lYpVdP9LUasQEc0mkPDzHMDScrrR3gA97f7lidek57BY9c4kyrHV9LO23N6BlJsyiwZ
hnu9vkpEJ5DM6fr2wMZ/sD3TyXzcVHR9eQ9uGpW9cDhee0437HL0X93sQQx3UTa8MUsyculGRj6g
8FKYlDQwPfZp3kanFCjr8gMje/g8LQnm6z3pyLq+gznmIlE5NXi0hFYnbOLhRepbc/ni5kR/unMy
sjKS1SFegqmQoTbvmwDp+Zz5/Nr6ihG3Muz8h+y92Ld15e8D2I1U+4bRo8+HzmWAsC4/T2u/BxsR
T0PvauoG0IeDAReg46339GC56s9Z5ZLNYr4xOPqedROpC7mEl35St2u8aXoLMaCU0HsUspwsX6rI
V1erDduvNzG0QELKs9pFp5gSbYa1Zr3hzrGX1+NBuLm2X5YL/4lQ4zYCwoz3UlpQy1oMennSYs9S
a8Vw5ANxBnFeJXRf3FGMAdhQObsNTaI/w7Z7TJuHEa5ffzmX5RazEiBzShr5VMSrSrbjJf6fFsTO
W02vGz65y+gFdHYbVIKY6d/+u32csDc29ryqDsdzMQJxENTwICucdckTxel1W9XuCgqcTgGa6BBv
ZT2ekuRHI9wM7JhLxdPQwbZSErcl2ipSHsKczNEoQADzt1sq68oeKgZZHq3Ddp0CVWeOryBynuBN
H+p/GGm6/lD6kzQcydn0dlTOTsm9UyBqdpN3MnFSR3Qzz75Q177SEZsdqh71YE79s2Q1/yvfJbSX
D4RoYBpgfUvODwE53DwMjcwsR4BqBfM46u9d2l+oaDenObgN4pF28OLbjgF4mayPJBlFgXrx0z1r
mQze621DaWNT7ive04tCbhRITO5zYBReWipnXiYk3FsTWeKc3Wgy5NjvaKx6koX3xUh/klaPuYn1
CEfxRXLL6BbidqsGXI6SLhOh+j1c3lZiPwhkqpwre9Iow+/KbnXNIfNaMx3KS/SXuHob16D0dT/6
S1OyWNo5ZXCXyHUgKGNGiTzI3yQm2a0lFZ2DE0rfIzHcQjuwsQbhGpZ3eZWjbE+yGAgtA9AyJVSZ
HeuwlLcAw3ixvLNKbV6CZ3eQVs1DswgXHH/J5/iY57o1tEkcFhAuoDNC8bFNfxKLiE63PvjMwrUJ
91GFmooMh8YmtI+jqXtZaJk0RxBkj1RpJ23ZBPlbQbcsXycdcivu2Eh8T2OnqY4duiO5PRsXOKyI
lb15e+RrJhHyYKbN9lfuqzxJPk0srZdPTGamzF1QkQVHAow+Zosv7rcGIyqzXxeYGx1f+G3Rs30x
CIuMeSpcWkbL1270TcRmdSRufeMT1BVZQIl++ax4jMvjF+arnmN94gC6joC+u/Xn9V6sCdQwtqnf
7bkE37Gf6eSvVNx3N8OPPPSc/Hr1gJzzlOUXWKC2kw6uUfYrx+ocRl+5QQJ9KRV+NMjWNjO8ZDUi
VZrxbvJeeSPrCObz8HVTahXzSvRbm3w4+iMfb3FLXWs5nkdkSt4dPltk2cQkMjHLUajFx9ckFaSw
AR0Nfd/1NnYYzi8nzxBcOV1iLoxl2IDcK/TH4Y4GCD90CzEgfd21rpwSthbDGsD1CXgiT67aPSWl
eWFewAn1y6rLvhjShLIyWg9ZnOK319oHXsVB/wfifLHgwFYSOXa3GtwRV7zKBuw4uqWmIAskNnjG
HBmuMYn5u3+gr96OlVZNmZCRGFPUyVgbrksgFxXqznSCL87icyC2pBo1kgD46TQgGifbtzRYLQCU
1P+52PGPxavnRPlPsnpORznttr7/fdEaTZn1aequxBycQHT1laVBeTwM08c2PzZicNCobeB3xd3D
2mZgNTDoaYzfTm4SgwxCWuVZSozh0gSTWBnXXPwveGr7Ig5kmsFKL9hJRqOqsqvvYtKxSamKBMp3
NrRAWl5sllcYyL2wenaPo+3d+k3CDlXuxThxUdRWfUU2iYcUkO6aIaH19wwJaF5TOkOLZqowm59R
3oTuNEYD4+777LKAEw/P5WAE0Qk6/di8u9CtUxg0b/YqTRZygHsxzsLZmo2UElQIOSrGumRIzUtq
zTQIDRJJH8T/gGWERjooFia3+hTYZ/3qTZoeLWQVWNuFDr98tbHqwDhn48EHcKHFVxlakRX5+p3s
OGiSOGbKkZpHGkCqpg6z+CuXwsSf3cDVWzu0SxVENc8ac8qas6Y7XH8B7c/7v4VXqqCLiR6383xP
D49/v0ay13UvtgribOre/jrpXIdupwtlzMkWoLNjGIOZeLnIOpEhDLQ9OeW9QMcQfK888+yJy014
EkZdkANkaVtkrziNJQzilURnTiPrIdYcZR+lDDjF1uiCTuHkjf+U7BQSZ8itOC+g580Ae/AC5RUg
6VUHNf+kccO8M+nuic+ap16LdycALtDdTpRrk4KeCqCdeF82s1b0f0IjWHXuOrRcpba07jQnBMP7
7XOsdITA+8jgYVoBruRp9XBjH38B0VVZEjpaWwbxX23GCIefUKZz/2FAc/TfVX7ZPqYvGi9WuHbE
orDPcokAbNCpWZgoCk508IDYln0NJANhEGRFZxyEBeh/aCaSEGx2AXJqcTiyrQ0/bOdlEThnJzCF
OKYH2woEsk2guwpNY5VGnwBw1HqYRjyrgwiIlqB0BFvw7Xh88oSVWs+itgjrNCOZZSlSbjI900Dq
MRNie1E3/J+oNgaKviHiq0niDxybwuu9uMFA5ag7RhqErDuwqONLNS19ZO0EVrcuinaocW1ukjl8
g3IuvWtgKOyybEMF+53VbGksmtlD6yMiLIVjYAw+goRt6uYL/Hzh6pF4Q/QekW2X58v9repcdSHy
f2w7CVDgLrCn5mDDIurRO1zDqsZWh00ydrkrV3eWzFGXdq2YVnOy6ZXUfi6kAaC3R/Hrrc2v0/lX
aUA9IS94UQWftnNKKZDB/xyitNq1suylrwOAwOZRzwKRGugS9cP93X/4qkDwyY/w+nEcD2t/KTTM
QoyTl1hx8BcupXlbGjXuV5UdUS+Jm5X7ntmLQuyzdkja8ainAHkvCLgvDdneaeOzsglpHNoh3A/L
nyueOHmuTUqL8kNLP4goYx5G9XKhdMqM2YVjSCv/RN36uImsWZlx4Kw+mCtGFmQDbRjA4PhPNwPp
2fgbUbXtQke2XPedt4DEe50MXL+pxw6HGVtAQa/OA2gLOOlwwvrO6SSn/ha9yBAsAKPaxD30K9jM
UQ5Euq+JmqhbhWVbTRUBJohHZZgkOHRORthGRb9CJTiFngstVdX+7C/1tTwEXwGWuMcdH0k58H6V
GV3e13VFEX5eue8kO6N5azdItl/AZJPk5wRg5K+OzgldNuTZB1TYyhMTW73ej1lM2awWiwHg0l4U
jn/PX54B/wjhf7U08eP7/OwF70FrnJNDFRat+rzkM3afjuFE5fboTpwI4LkRA0/45oV7tXP2wgR4
rdk9lC448Rr9LQzkr6Ei+FNXdNtbJQrZs7xO/rzpBjkc1jFzkFeE8X6RNdqu80anLTQlfxj3MfXz
8sPxVjd7Bvn0JW4z/STJ/xFlZx9lKSRblUEEpD9+lA2RLdqB2dBdW9C/khbVse3Z6Huknnef7hui
DcdUSgQHhDafmETK4TJEGFRfuRB7eRWI6gMHJbL8Yvbx/VsS6MalgDm7uMtzyoP2qzgpyTje7g69
YlLbRF3h34E7Ejj/eVzwgqAOV+vUSG5LKM/gN2Dr2Fa82Q9jCOJgkUOi4z6rgOwF8UcZcGzywhxJ
vnSuR/RMw3vDHQQMs4Chcj+K5oL/M/QdKSle9D6R05wNqMw66B/iwrmZf9TVc7lq5Pyxq7dAktaA
gF4x5EYV9jOGctaW928I/AVRm42DhrDBWCTj3gho1uejjbPrumbIHexsUqKPzGAccwPsWDVXmel8
dqov5agedhljB79odFIIXUe6eLYcQtB8bFyRgN141ztuu0Nw7SR3ecCOf4ReOnpAddPjZl2FXrzw
EKHL+4PRccOfaEQO9U7U6//Cof+gWdQsBNx6tFOOgZP6xCER5fqK6OY8vUGhRJ7EwoOqFM8lYPAX
U5XIihN4Nz0Ya1rsd8LW3rlo9F8lc1WWCo17bRHvDUB7OxYo0S9JYwQ+G/9NrqD5zUPv4nu134E6
UJGUdFlLIFYuurWDoojBDzzpOWnqzdxrZFDa895oDbVT1TfRn3PMDth/YRUNNH7jGneATmgfl+AX
B/oEinruovOJVTUg/ZdhMcYrHwREJVkXkZgDo03hA6yHpIlXmtVWkdGnbQDxRS7+ufTVnUQsjxIq
ZT72tDpATOphQgSq5Wl7QRm9e1Pl2gg8FGkK1HqXEn/Id9diV0CuA/rl4LzbvtjQ+7lRNsFEytYN
IGU+YZ2FjBaQp7HR0j/Aizh7e8FVgaNtCoQTLWD/FZLKojUKn1IOM7cOd3TgxM7mhWHAhBt8DPgZ
ja8ALwdCnHpDxNB2VHTa5aI++TF5qrpA3jd5n5xMwxvITF5TlQmZ7IBQEAzFqa6glCadYQME4VTB
raBEu9RQqRHz5CUd2C9xfbHwHujoWdggwvc0xjDsPcRWciJSVovycfLB0wa+A1aMHGYbEo1+7tFn
1A8z0Mg7pyTYUiFVGC0sCPsgxPEeW8k5jILwThAdL9T268u+eIFGfSsq5zPYGyS8+mmaeDlgp+LU
AyidwH9nUhCs1+lwvttbdFFc2lO/3sFqGz6z4iGqCRMAmfDlXFYLOO3cQJTkKoexXSsej2hQfbGu
88x/9R21X0vrfhjx80iy7mIsLKRROwI86lU60mArvGIpW2TJP5v+hsE7T2+k39ZN9FtqZ0+IMv/u
y+1Tv7adBfOGRiiTIGoJ8BXBkEizgOHBAvYpv6Bw/KMaLxG5vBQZGKzadSvxLA41wRhKL9t4J7UH
Sm1cWLPol2nZucjIZWPRs9OESCIHQPRP/prgHaBvTW1f+r0Xkor+nV4O+bIbFlQuAnEUmSek4r0K
ibKu20MSVJACXq1LviA/99NMElfbAqvKsn9UxJSBx3Zzgw0HBhyigc/ijCecDrgSpqGsh3ceKFie
rvCeNaJ3t0oDHfFoGpsqiCIdWsKjXrmvAsHGaBftslAJNYWSLUNQMOyEBt5bbAlx8lOWTMyu+9vV
xx7aMqpvz7FmcFCjClCryIWalvpwdK2UlCZylbRZ1LL8KJD3L3i3oCu/xzHEjNsYlhFD7ay/3jXL
6qNBjUZql9FeWUYPMnYtNvhIyP7IbeNzJu55hClzDauDp5+VgPmMEMX3GoPTP4kw4Outg0iBGEHO
SpyQKpaxZvUSW9JC5Z0UmTzuF5LWbyKTUH3y0iz9xT0BVzAjBQdxz32gdWMYqm7TpQoFq0iNWJr2
KYqnfYCDGegbb9ig/F9aBJeQ3zKCydT59+0RR/KHs1EadXY++WR/reNSXiR9eMXBA/YF8K7IlgC9
+ts9pRwisRNwuLrAXmZwgj34Dj+lae2ehIYSSKGrM5TKLgRIx6b+R5o+lavYDt4AbHyW+94+r/Lm
p2GWBmZEzvpN4UyPNpyFai8Uxa52yoP+H/gS4o3Rhbe+DWcExEDAh/J4F4DdzAh/qaPbLvnu0Baz
L8tGnNjnFjm0LYbl3Mide5MdrsTIEHUFi9uF8mb1HqUwEnZ3lZnFg7LXi4JvAJcumlKjBEPpAmwX
9S3WE9I8iIh1GhMLTx0OYGbPunf4UG0TJ2GGL6GXsAe6x1e95F7yzhY52BZJto6Ln+6uS/b1ORGy
UaaDr4xHVmuIc6x6hQ/qqPmxi8ra+4abAxcTrRWTVFG2HjQgIO8rBzo+7Rp9q1SzvH5QzhnEApK4
GgCILQ/y7H0pvaUCBMCdh1RTvZnX53DSOpQ5S86Uuok5bjoyB0jwFW3/ySpBgX6J/gJ2HfDg/C1/
uFS1awL9Q+k+SzX/CBXOG7EGOfpbsbxCslbgkMl4E/KbFPWl07r7CkB5qEjN4DM+12vOINMhsK42
UZp7RcX4CYrEA6tIh4keDiQ7+EsK7OKzOJ55QUy89JHZk3ku/HJqvbsDMDDmTd6NkYTgti2Xs2oC
b9dvC4XYsSKLJXrMGftOMF8T9ecogAbo2iekzr0PiqveqYEO1OcVpUkdT8n4RGMl4qFldIozCMy4
Vz2n/UGVc6ZcmOPXzxPtNIYIlG8RgKjUMIUhxvGe3zmoqo8beS3F1sZSNyuM26eavT8hmeePN5uP
BRz87CkNVJAjD6XDQIfzXVivAwV/3jzLJjisKM8QBo5BSpQPVZ8585nG8Uc1IuoOcUZmy8FFzdx7
v2WX7rCP0cQKgNokfcFi6OtH81mnffIn8/QbbXpxxMwLxunF9G/qf+wAbOHTMAsda1kpMQobATL1
jQR6Jp92ys3DqXWNYA5FcxCHNgjVmVTAoYZc+ayOj9msyl/VGmoYXlV9uBC4/dQsX7kcF9Xit89c
Xj1/KSFDPQy94eTmg4Cmcwdu19MbaK8uTjqz7XP9PTDnH1cOa1gd+TjhADhaDbJ3fW2SjBd+gbZx
P3UyzJayAQml6DQNahF5anQ6J8j5Rzm1Un3QuVxtCx6wRweffBhZ6hcTVSp1WlbaJoMFccn9w5oY
xn8szKYw7m6dmZI9LYz8HoYJ7fNzzfOR4V2GtzjgNyTEPZtTB0WIe7oww85/QGHJFJLDDnO1jtnu
tnE3qCgeSJfu84yjeRYjJWf5jBp/Pyg/3n26hYqm9GR3nS7+BAtorPwHQ74EsZ2oyL91oTn2Gr+H
o5LrsUnBlLkbGgEoNOwKBDq3XXC4faBDZvnRVgQkPdGlESn0qfp5svWj+uMPm6M7W3gy+Y6syBVm
npF68+TCKkTo4NoLhf53ICLN4eKu3ABLGCcR9hHWMZTjqPi+RohOGykHsyshAH3rO/XOugXfNoDF
Szn4igKlDnjPBLS3XhCICNE0l72b/jU5fvxroM1pP2aMGWBG9Mh5K/0g1RxdbO/jsg1031IcEDkv
CECpp8ImhhWGxp8JA5cIjMqmU4qpNfcywakboMS+Ue35iko/INrGEuabr/d+js9iqcUeyEXE+Bb/
pMIzOAeDfjebze/H1L0QcE9WmfeXLOgUAXbbGLIfcEXC3Do2llpi/sZ/AQ5WkE11vWNmbccmnb2H
n7RLmgvEk7H7Br1Bn0Dyj5BxM0pZW115lcDbS9aNdJGHvy88XFVJEAr4eVWCy5goaVcs0c345YFb
jPWIoytzeC1N606Cg0Asm8NrmHLnLjvDURaah/6HCJRzIOF1YLijYDxU8TAweeFpQfJRQGlh8NT7
czNrLiEgr9H4fr7qEbRuE5lNaIW4Ips4Lp9WMLn/nAZKaitpNlJ/fo3k2h9rnTss2NfgUP7s1hk3
eEBspzKGhCRC7b20TgRFVQaFlXUTleBEPAPkJr9u713LJg/GdU+oVQJUTwBwdWP7I6cB/7+syFBP
at81UuSn66bDbBJQIZDse92+xpqywgMVgrgc1wkhqAI8qZ4iOW077kfjZcRHdTiNENrfph1cVkNF
irn/DngTSMx84crsBFqFE63344QYKp5ty2qBjaODqRNuPlFDZ4/irXtOjWFDBQa2IM1t3Mxot52Y
BTy+EUXMRJVQbnvbEagVE65hvxWeifJiX3gGQCu6kOrWc/7vxTG0QHHftxFVS0JHA+vQjkN5k8Xh
NoUgkEXxN9SujLTKIEVbF35bpsXoQCWQBErpq7+tNPcyySeKdr/J7AkwjbUowVNalgYgqLfZ7oMI
AUzWoxzcwvJY6xCXgtVlwO7HykqqXOJ/9gcHe2Cs+3gJ49wBEPqgd/WMfpU+dsvEBNiBf+/Uniwg
+47VjbcD78xSfXiTjxdYKlssPxGDbn4Zh9z02UUa8rdM6pRjd4LICQBvIjps32K30mNSP73RUzcc
GnEw0wiEm7zLxdP73AcOkI6XCtiL2WC9zUuPPX5ffVMXeaLmsJ1p2oxEm2WqFkCLHGz8u4oLO6La
aw2jD0RaAUZQ1bG/OqM4yXuPuA/YIXbg6IaNnidHj10tW+YZp1kjVgRfo72pBqLvQcCmubLSWNEI
3fUeMGlDaIfuDeir2o+6PxTyCOQJ56DOUC0xm4cjHSy5kQ1yszMqG6i8ImyGTUi9SrPdnNz1uoF6
Hv8pCA+rIFeXXz9lJLej8DVc+Yf/HvExUG+xCeO84QguKoHrbZxBJ7MVrNM3AqXG30msEi5cjX1t
92c6auITfgn/lDO+UNNqeOq9amZH3TufMLykbC+JNTmrc7YQiJ//XiYP5+I5CVCptFzanKQ2BPsW
n8Gb5vsLGsnsWj1b16Vjfp6EaGTQ0T4hT23mz583gvIAXjc2hJlfKxNVkPTEOenCRtvIm01uu7ga
SlFitjAxJkny/YfTFQQYaWGT3uZjKn5vBAFU6LKSFRn0sLxE3zu4y0SauNABQwv7cHlXfDyx4vyN
IzrExytp30pC9nBpb04ur4Fe2tRKplIzdK0Ia9grOLw3XT7RonJXEBSuQ7wDusdsd82V8220GXyi
NMwQdnFICNYvWC50MVl3FC+8HJnUjJHjWc1xUmlDolp8I+OE2NgjV8vtmgzUNdYJAkVjjhcBFpdE
YrYTvpucjnjhZ638cGMhOLmHQYUVEtBoAX/pxLSxMkjwdz0SDcgpW5p4dbBHpgHIlBT3Keyw8f+I
nao2bgs4EbpkUIZ5Yic0jHyC88w2e+Q9/yZI52f9AgEWPJWm0SZv/iPhJB5OcmMtOT3cBlLb1uB8
dhDl3iXHmFMNIcLsLl3qHYG6Uqn6fSG82agCuhD9Q+xEaOK4wshu9+EQOLH+F7DCKREqMCYy6YWX
2n3bKMRFpmiQhhpCe/ZJ8AK8nq+alXmQ2jngXi2vrfZJxxaoP6WznK6Z1VFnD+bDluk825Xxp2mV
51drzrB7+2NYoaAl5jG5ugyE0h6DdVA42ju5MABxlAZKarUUKiyguyqbKeqZpd/VbyZv1WHXDFzl
tI3PvA0WA8fymodKfgqpqk/UhHS34HxWgLMHjLCoHgKayYyL1zQCKdiFzKqRzNUv381fOQh6FRag
DMy7FXabrxXU5vu4tS/BRX2fdE3oaeGLtKbeeXuW/xmh8u5Zc6tswqCyqprtrWjkc89BRjfjNG7G
7ZyUxtVFm3cpZYknL7VoMlQZqASEcgf4vKLBeXn2llGfCom7SFr/zXXSXRpQczMQvSdcrsWbPZgW
G6ULUl4/yhzPM2MwvP6HP4ov6k41YH6Dof6G1Tvwf/A3vdKFfFGdSFpHVOyS3ME9AzPhr/hi8eYv
8NcqnciiMwiuTaNgRsFSaqVsw5dLMv0Nm+vyqZM3BioqL4ov6zrF8aWqfxrBbuyhIj72LWimvV58
J93YtjEPl/DyNfJjNJ6VIKCN6LLG6NB1+U6oX9CkGXi7P9PVe8ITpDEvGlKYefsw0iSlbVzdk4BU
HsfBGUG+TO9rKxRlkhAp/GYO0WXu8ZgnDBNSjbxCpKyO1ieL0BR1OOjf/YlnomRowZJrVzrfvaPL
X0bKJszpywmppIy0pcDdKduP264XjF2WYE6vOt850us5AYkOgtm9Uu+LL5GySVfqsh2mATHH6Epi
SiDmlnSEXxg6XLwmEWHb40URbDNzxlfalZPiFEjucm82LrSh30IzOd02gnxBDFxHSid1PCPkuL1g
F8aGj+G1fklGMXNkc6g86PjzkqofwBJTzC/RrHAwXgzMXxeO5PTZBltMQIJ/KyalBl503h7ffdrm
xYK8LuWcTi+ctSxc42Ol7NgNOuaOEXYb/LA9Ka00k4jsvrW7DKiOHheNr68oI+7y9avVwaoBVspV
6+b3hKdE5HtpoanZBCBlhB9k5DwvvcwQitg18FdT2/XcrPZrneqCKZiy8XE6of28quHY/JZbOqWE
DJu9jh2BTtl3GH05UX8335CaAfsQiWBCHK2ifjQwDWD+5H2Hh5Xu5RgIsilCCC9laGqVbBFpbAlv
OQ+iNcRE+3ibrQ919eAmkbEJik/p/7xUWcFCsP82b+YdTpit0rsT3E4xireWRri4eMnrgpbtHEbL
shjq50nsITGynsapu5L+HzxXnjhAjw7ndUapXba1KXKTgAupk8WDWztE1QsqujSVSxhrq8qUeaqo
gSlS+4TncmxUvMg26Mf31rCAbuG692sSawsSDWviFXyezA1HraezKIjW2FYv/1Rp9rxgEV9odl1e
pfVmJOTo3gFJDfrS16ik7Ok7I7/FjB0WjOUFCmNYk/fWcQy4WFg7iILpWBUshrOuezrx18Fv+9AJ
cpjroSlmt1zjkB9YSXr3jQWVKiTq9C4N27dgPTfATBuF/hgMHFT+/R2u7QCpN2mfQD6X/5+gVURe
VMfOAb++PUXBOJcj0Pfwc5GJ2VwI2M5nH69RLv3mpNnW7OySNHDfjcFJ5PX64X/JJFLxsgV1Y8t1
wTNUg527SdZv/NOpyOWmbVttaRRb9kpR8CvcTXDRM8lRxOMz6Yx9Sm/bQz3+T5lHp1WmMfs1UnVS
wu1+ac5RSK9n6XDZTfamKCjzJTbVivq7VsYVr6Us/InhvR5ppBWju92aFniLQRIUWUDJZ5vdlZPy
OUH899mcQpmVav+xveoSSURH2EMvDybbE9aoSHy2VIiPsftC+/yWgEBLBY2Q0V/7AmG6FcfK5Quw
50pukLvucmK6V/HZ190DU1eHIPTHGwdmGv3vN0c4xdmHqjpIO2slrZnPGFRZDSM9cK7Kx8AmUG29
z42d/PSvjafk6QRYaQYvHgb8mHORu1ghfPSve2/EGwO0ZN+qcQWIzknk4VvbK0/8NU17Mr/6io1F
0Lktufii54MLGMB6KpNPcm3COqibQJR4y2gFMeDLJYe+pS0vwOHTcZX9W6IdDVYa7uCTsNxwE/PN
FH4O5kY+MMs1j6PbgVUi4/4/tS7m7x2Qf1+2jSpxTvhNO0xZK6MXQTycOWGbq7QBggQrrZB2lS9p
WnCZY89RYa3SpIwQ1mCtcPKFyJGJjBv2yVTMeknRx+oPi7ef//2GOBaPjpSty+0cSN7wOw9l5F2v
dufKn04cEsrqjDWoUBj9q1ZlIyMBzjZs73rDTNEkfqv51VvmYl2NGPcPxGcR738/M9ZDvmlf654a
EiLXXDANMvlzW0fxme9+3zC0+/DWDmLSesMwyEHyBiJo0ACYLPvC2DjZtsTaNmyEoXbXWiFV6udS
RWAQOtKXtAXOEPae0iQOhZR5ABaIBoWXN9PHu1uj58ImC3M15ADSemb4d8kOgw4itblYFCL6vuV6
XoMJd0Z7+UURpIlK6k3rN68d/GIeNINdPlw1Jbl+y3KrolpNCdXDZM/uoE3Nm2tS+s7o7LDwpQHp
sD8YukWWrm46Xrgi/6sObenlEYosm+pJr07FCB4EZIwC/0cIMVO7vk/nh+elG1ksh6SfrL4boEcC
b4ibTFA+yMSQ9hyAkDDNyuH9g5ymidk5hpze2k8bP0Uh4KdSN57k4DlwDz+QuLd/BCmy79V3CpyJ
9zt7aRf8G+DMZdRoEomy/pR8NNaEgRWuUwt0TdYdIM0xwy2O18r0TM8MkxHQ+CS4dWeEROlVsyFc
Hr6zR27Bzd096taebqSaBf6XtnwKwoUm4bUGapkg0AXIzU0GfDfHeylKvTqYqo7ugcnN3WQ7r+l0
C57EJkYYkOF3yj9TKANknRX/fVRpGHtf/PYrlCw8YDbucAkeyBdKmLXsBHyNU6Rs+6gsUg5+ubGv
K2JRHSu7xtP1V5AmqMYFR5n6WmdQux6oYtlRlt2SCHy5dLHKnPRgbBONCKIYZP2QqBHsQADTUZNn
Gj6xqC8gjZnAQntaichd3X3cDDYjpgchyj5sRBc6jbbhgAdp44hy+UTFUCobt7zRbexp66aN65py
d4aMJNfF+MDw2AI0vgI5P6nLh69xmlkROIHjUT0q5J6AdG7ghgtNaqRoC4VHjcbVn4NXPDBN0PSH
ym8M7yNSxdMzhdgUdLfLMpvP6n4FIck7Lu1BfDX7dTI5y1oiaJaGaLPeQnThPNA/b9v7Ky2ty18U
zJRz4qI/Tpze4mJV9ylwhfkSriK1UTE7cfvnqQm4Aw2EhI0o6vyHjTZGzM2RsfRvZvH8zIAfshlW
PvSF939lzAfAziiJ0QHXZtna+cI8iGmVOBxGES0X2QAZJS/0KVYE+vzg/UtWVL+hCM0m3jpmuHct
VQNHAIPVsmtjH3lZ6+2D0IQa86Dr1FVZvzqYenvLHiQbUUWjW+EaQB2h3tUtmte3C/nqmELG75ID
VFqLjCiL9XHx4UzgZC766WxOUdeRnfywJx43OFptfwGiIXNO4VMv4cn5bEmaCVLyAL0NlmZlnOSp
SjYH1t/4Gfmpl9OGbw5Sx+/nrgdMoFuXsLeBTyM8PeiGT7asNzafo8PmopXRFRGk1k8tDE9oIYzS
RiFRTnbdULYEtxBHx6QOwv6opU3RDbvCKNrgMizzOhOsKCr2GPghHiokhZtHiGro6tFD1916Z1E/
MGilEBnDbg9+Edx9nMhYPv7iurp6XSgfVG/7W7laO94KeA0YxkmfJwhqtBPU3B5UDcBOjDD98SN2
ZeLLv3XZmEOMc52tzhb0He90gOf/tr30DzBdVb683elng9+73pPFgHd5su49PG5i8E6N96Wqmo2J
tPxwvIR3BoFdBpQvXAmKe40RNHLOrE3uf14A/QSIpvgQIF/9BN8vu68hGsxdBiCRNFTxTGHx7nTn
TJ5t/8QHO8UNpd4RMZRJk+BlbnY0zzSWB+wfFBX4I42f2MCLdj3xXokmhSqImn3fZ6mUX5kHQVYW
YkNe8MrSr5R87loePUy+4XmyDbJ4ShD+A4/vf37mpnJksJZeAThD1ouX5hR7EV74rrAw1xOJLTFF
4RNvB3ITZpxjglmOgiykX//MggzE0yvcLe7ULzM1dEJN62JQQHX4hDtZM/S6wLCmi3pIAcXYsfgH
F0gEHwm9YHIaJLzHFKbz2dlmq2fl3vOpTRoQAnGXa7/jn8BmRRygK79Ij7bQjLTUbCuryrcdszw/
OOqu/9NayKTj5BTUbF0X7R26442NHpHUs8650TNPXO1sfevTcQizD3fHxpgofuUf+ok395B4Wp7Q
7ma7eSRst6cegqPtIaxXplP2GsKqoRTl3WaxYMtyk0tWqbtsJ/5tIes3vR/GF4HvYkUGZEF+AHQV
g1Dgn5+DCUsQkOFrma3d95DKux4SiZEohpQ8nMLsdbbuClBl2abYFuuBqDrYrhGPcopYCUx+UMSM
Wj5vnwi4VO/YjlJh6IVxoJtRArZYfpalQbbUCDJswsn34RusPNDe8hSqpId8+5LJhqA8r2KOe9oL
iIKkY47QymYVUgCTqRdWWRCILP7IqoSVmXC7pjhqIr/o+YuJK9iji827Zg6teXOVP87zCt3TCi6J
hktGQzMo3UuuWUlLYCcs6rvWGb5yEYn0gVy2onewH/LnHa9jGdFvDTuM/qWQxLzOwieQzYPz5IR8
fpDKiZ7w2z2Z7NRX4FbVauf/99mHnf4VussyikgPLNJMSYhh4334OLOhjsEZa981furitTRyGWG0
hSCWE+Fs0grgu9HVjdjY94IlkUr/K9cRjp5lvKSV+T4XwMS298ReuTOgsADXPSKgMxU5KvSquREH
LibIZLWyznGex5Kon+imkNfl3BXYX8vHvh72WiIm7QQN0VVHEcPJ+o9lxrOnXK6/NP4uqfdK3yhs
gCtkbvN6+OS6N2pPUhrPKKAevABGcIEVedBLH+R1GaBRp/5ZLNobBxRHA1ueZYGL+PDnP+LNnZzL
xy89mfUDCG7sZPEEcs4qPzP/QcGvRXuOqKc0L420PRVMwT2W4VF6Fyubs5RXe7v7J+RilUoMP/lY
No1RULVds0W6TESTIkG4Dx5Ff9mFnRPhWk4Y6V/K22b9lde/cfjDFAz8GuwS5a1vwEvUU+YTBBMl
XGlyKtOVj/J8AG0I8HD8Kprnb9ZgtU/R3379fveALIbcEy8wCzV2lD/Qle2dcFijXfHJB0OuE+Ni
NLrINhYXqMFoCx6TMEZLRSCMxGOl5LT/wmNvIDEaf3YJnCTNn5bEQXctB4HYcGcohkq/YKMIoq+8
/8/5yMDEbxQjw24CjBoFsnNMdrmrO6b/0QviY0niMMehvjs8yOrR8PrnN5reyicVS3Njzh0fsCZL
I9DjxCHsApQyl6vZk5xNuwOSjCSxZLpOKXRn7oiqxNDXLOjuzCBKAo+nWUur5s5onMQFAsomQN33
G4jBkkpvljQvh/hVi6CK9I5CFUpm5gWlpv7peDkvxLEr0oxyxZwboYus9VWLEd4Q5qE2ryDAMBmh
D0T54yN6blAeE2ry3ruZqiIuDsbLR4czyqljj4G+dkm3/03ZbNFMBkPU7KWu7ckXSr7zZbIoJjHz
pvqnBQXEmQMxTonfMjehexqfLJGq2eBofLb5PMc3by5VdggQZcqvgXo6Nq+bQUPAqquKm88phWy1
ePVcHdIoXw+bWQED2iUXAA2BoW+nS8S5YLutDcOSzXGDsQUklU6NrB2ttijmgpWHP+B1uHvf1UNd
ZOL4/LhRluxITZQAeIhbyX/zRebrzJoqQlS1Qar4tJACl7YT+BkGFOehuHzSvJLxS5KeYNu19tuk
GVvhHqR9NR4ntsnQg4TFK5sbX/iAcjacWPO9wYdtyAu/RByhqSMR32dsELsnFoxIhXuwyZ2P+Zvb
S8sq6RRfguMG3WTZsRigMrOvabL9+WFwBo1MOfvst7IL7lc1X+CwQAB5RLmKEbHs3DN//dC1Wgmz
W8rs24Ok6htJCDKCyeDU6+NmxclmoIpGTgIpoNsVpKGyHrmpV+klAWv2ypPE2ILrQyz6+wmrg5ch
qwr43wkWECkhJmwjgPqMlkz8Gyt/WvXMC2GVRwcPiGaP+RG7d6PBq8YccQ12DobFlEKkYvnWWgVU
PepHOLhI53OHIOHVfVKAku3KRCQqB8laIKb/IZddXf/q2DJAi8coMn9FfBuXAcnkw4e8G4knSeMF
hYxSU2kXmeekf789Em1MpoH9u6+jjo9tZM5URl7ioDVRZxRIoI/iHVJQRud1yGBP78FK/PfQFw89
+WeHEQ/ZcwUS9XPIU0Me7t1B9ndk1fJAM7sC6nGsDA2QWL7YW7eHEPMzrZU/WE3gFpHoPA0OJguE
jICv/FaJ7b1my6UFQSzEhh66mfUkrP8CPw2SRHaTu4HkPJWsM1w0K44rOEowjg6rw2L6nz7lt8N3
j+/SL73RNk3Q4YFU1A7H17BEfbjGigs65iFYVSKiBiuffJw28JIU3wqFc3V9n+4n4gAL8/XCQMF9
QK0Y0KhuJ0Jlz1sXYSUldtPcz24POm9fOEeHjSvKOgAjxrRP6ifl0//lic+PSLLVtpobEPJ0dMnZ
O53ELxurN9L+tSZ3fVGJagHNBIMCXSS+o2HkRWAf0ZyvitzX1JP9dBuf5CL2h1qAIg3TolIFJ/tj
rsyqS1VxeBBfHkhy+Q/8Nm43DYSy63YTKKCx4FLUMpCsgxN6eoHERqfYeL2RAWXVsqF1QB0/6Mnz
XIa1mtgsgoEidVo0KZ2FAUPk5lcFakl/6Ruw8IMdrjCEz/2j3jt0qsTM35TSUhJBzOTSVKE6aCGb
ni17g9aKP/ighYnRTAW2dPisGNezpt8sXF4YEl2pBBFBv3dxmY39U1+w1ZsgCqrCaNV/zSRu+nJC
oO0SQ3KSxJuzOw5XPVgvdRn9Sq0DbBkYUqBFhCfISUFhXp4Tzo1VrmMGQIUUk+3A/7SklX5bSunu
IHzjD68yz9IkWe8LZKydkeKwo2r/NT6i5dwFUp17pYdzIAPEXU30sQwHpyvodxW9YbZQdqAM6Dfg
BYLiSTaY9iOqdqJUMY2Nc1xaiOx9POMkG6HT54QewxMrxOUv+QesBp8fmm25+7ieIcn+VmdqyFI2
4bKHZC9j/rpuN+5dBRtvL5CdM1q6K2UJkXC7cCBl/EwbAMRuRIMMwMtWX0WsMxH0+cz3AlMscYt5
kxOKi4GAW3tfgtNw/FKNodKz3rZiLphJWZd/9C9xzOGBVfyqTeRRC3Vqjs/Wl4wTVHDJzs99BXIw
oniVVgOkKl0Ino/o/D2ZAoc797zKggbYywTT7I6WM8VwS2BsAtliZj6vXuEKXAEC3Zmp8hgGGpYD
sbeMvEdWJuTKlpyBwsXJt09oMiCSPfW5oXS722TcrHhE7K7hhz+ejbAILzYMl86IyV3gXhw5ETJT
XLr/uDPPkv1qOfoQJw2Ca2CWnhY8sXxfEpZHlMJLaZ2/jac0Vh/8Fa9bZD7XhMQGY8I41XcxbmE7
w2XtFhq7f1KT4iIQs0pcfKohqNYuc6fRAiulJQxyQoNEESMSDffuAgwDUqOOLLZ3UZhNhShLrB2E
3xcoebtYgYLFzH9vvexaCXGQFd/Aq3W//WCYtrSj8l7QIJDuiGlhVB7mW2bb5PjWTZyuEPqxmNRs
lkTZmAg5okPZ9KLV7tSPJN6iZXgogJ36u2vQmXgx3RBqlVa9TZ5Wwik9uBA2ayfZ64BBig31ju3b
NYE3FsaVVVM5nIuOjZO6QnDpD6GqBb8kIR+rvEWXFlwWYEOQZvA4HjtrAcp7ioa34WXO6CXc5AZN
gWfKpjpX/EJ+B7EmJr8Ch++KNTIpo1hRRMc/PdqmQT0FmPu+0vFJMYUyC0ypr4piExMVKIhme6J4
dKCz0w5w5TX+Glcqxu7OPdJRQ+srvKvD8xFBIpN4NsZnes7cU/r2DEI3VkBDLt/x7icm/WAriIyJ
iKnQe1iMfCad8RWcuwL6pAQkTlVahlEmWWTBQpY7BNh/J7JM9OIg87eErQnmSpR+Ftoc1ohFx47R
tG/JvS42xLanSb94kOFlyR4qosuLdbwjD+l5SVaf1uAPCoKkyZtGgVfD1/CC82aZA/RclWxGPrKz
/lw1Wia4cGUmB+Ry/7pNgQ6pAlkdc1KUpYwNLkCKCWvDKaOOHPpBWCHSDCBl77Kp+zV+Splh+Y/j
TiivMD6GKXAK/85Jo+HvkSb+dL0RHs+eJ/bXNVp3m3qnc1Uuj31odnhqh/H6y/yvmV6QWAOlEfH7
yaCuQzvD1fcPUr4lPyT+mb3NPCKI+GnjZzs3J+jyCd2qQ/z2xNzaSH+KQUFNl4b387guvLOBWqWu
QBLsoFaXU2VXIYt0Wo4QmNZuTi3nyeRakykahCRVWKaoefJhzx9GodLU8wFFAxvyyTvMTM4JtPB6
U5PZQBl91KVhmwEby2FgmZmZNt9Bb8JLgnpIlw5ilumaz+VbROMzFgce2dqPHmnWxj8gIOkv6xWC
giEfXzK5CspgwI/tvVo30R/jxSIRSDBwmRJOOTU1shE2jEqSt8j9++FsXVP0PgxzPkd3idYLrOcP
+Eb2LzjokjLvRZnR4EV2WnSy5Ybfh21F3+aF+j7k92AS/vAYfnSz+6EBjFwpJyfffU5MsmGWmLhD
AhpPZVXhLZP/2mja/2VeHLo5MlIHcqxKu71AIx7OBx8pv0lSC7/Y15jpT5gVKa92BTAZv/mzysuN
0TbpDm9096MV0OJuh0HCKfJT3OYYhLVx2MM+Z2744AT0TN1ir1J89gax9cc5ArygGeu8yIfE+fhO
ocvODtCccPC539BttBt+YVOdc43AzhRk7b0Yot+RjVi0U90c4UjJAf7kCI+XzyhCcC5P61Merr9o
yq4igM4VC6LNVYWeoraoeUegiWGLCcNbzHVLHpsixGIinfd/eufbZqv+sFo61pX/E0m88jJvyNlK
4NqnZptKJ3xtHp3QkTjxwCROrdc96Ot+LWWkYkJEY/JmtDwONvRVxFkB+HbibUuB035eRUaQDAjj
85d3KKsVsyqvRi0PMYW+7aO/2/0vvHt6F+4+kNZEnAimcWyulLYfAh1NJKwRdGvm73PKQO2a0783
o1lFsXUn805CcygfdxSGAb3gp0Iks5kSw16m8DiJ2QcRxIs6LGTMaAj5nPX35iWurv9dlWbjv2I0
IroP4KLrFSIew/aE+WtoKmljm94pCswurvccrWfmf8AkHwOrNTq3hsBV1U6bqLxNmdBtktFDUpMr
IdPHhLnIQcEV9wA7g/wCa20YXTwynLTmUODq2LS/tAvfVEe/odcrHxXISGFZGycNOtusQNRaKkoY
F/Kp2KTPsCu0KTX5fXkb97nELg70Rw3aho75xZUvEB3pjyzcMZy7Us6Iet4CMDWVx6yzA9TGFc/g
BD4XgWQ9whDDMWPTjXPrzbeGY6jVg+104lN9DYRX0a4fDr7gERRSSXuTPIImeMcwALTnuqVwE8qe
1rKDLfFiBx4MySkb2Y2iBqtJgjExxo9xoPhANj7Ow0hcMpyVRrESjKrSIChDPbx6Zm0aJ2xAApuZ
r0tf4RrQJxYBCs44ww1KG4+T/H2oUka+L3i6y/s98rB6xQPTV1KbITrUfUcWYIMugV3AAbyI5Fkk
/e77j3q9gNmA2SSeAF5SeuP2X7DJwMY+KJhyU9NDYbl1rbOwjjnj8mEixeP7uucxZn4bAL3FfNR1
dD5IOTr5tX36/ZgB9lDZI5iMmdqN+iJyNpY9PwUJ5MBQoh0lLtVX9o3HBv9Vb47lqz0ZBtykeMFK
CezvDUTi2cws1TZBc5q+nBIIyKIFJDQt+B7E672aLceOaw1G4MQJc08Yr3Wc8HyPh7oyLLC9nvNa
NKfCl48/GVKObp5V4muVuj7KTgKtiCH8L5Kp4qSyIYBkySUcDF0DwvEVS0hJfkD0QLJS7ZKiKreu
FqxSiqtpe0mabislM3JMbylMXZQ4wFQk2v+xueGmS8AvIMGPSVphdoycLTtv/ouE55JVY8z1QxqE
D87FAWz9OUg4W1YfmRH/umEh9wSIhdt//yQQkODbmVFKStlDdS3XlzH82ym/feCi2gc0qUBknM6e
5X/OWty+dj0PygVTdeCSLuDn8Hb+hE0Il+m4JLjEJzYQh8/pVnfeQSwYaTnPD8U1A5BhMXIo3JM2
jftgc7B0NxgqfGVNrBKuSkJZ5+o4PYcQIehqLYWgxfa6iXxtXhw+U9AkirPJGnw7cCSnOkEK6Vx4
QYeafYqciMl0rfLK0FGGVqTE6Bs7PnjeyIxPguYANBQV/TtKj3edBRsHeOli6eeKmtvxZ/YzrW4N
+MYeqsfb0Crsz8HtmFhh5oBEbRKll3WceT947hebKYmbz5NRJGeVlnqtCO/+k4454umwQ0zqyF7d
l5eYBPqWkTMF5S1QUItlbcHPpMA8c0sneiwomnkCPOwFbaKM8i+oBT2ikNh0YEXdijMhn1+etnhj
X09+dbbNdbTxaegGgh7aE8mgv8umv5NWYOcEHfcT0zlwIH9w01qi96Z0DLkaXEiQ2myVyVIFbFf0
kg3FdRc2G369RZGgmyPwV+0l8/3l2OendRuJbWwQ45HoQMCYPPgla/HcwES4j/SmslONNZQ4ERuO
72oHe9piFT0bOIes6gteLWoFtn6LS+T0EWwyhnvraO3j+7fdUZtCzSC/Aq5Cr2K8A9I/X+noYW0a
Y72N5R8Wj79ipH8KpnmaHk7+DUP6hM1KXVnBY2+hi4pw+AA0A3djD+0SIHYJ4mp/fO+FYKSWzzAX
u5MOd7LQz4KQUXoYWVCdEyRIR85yE0f35UnXA3kzqlYlOIp5wz5fqzV6HvL3X/4SNYx7Avwzkzhi
kitypgJR/h8aO7e3QSEmaYLuV6DCJEIMNWE6cBisUW8dkfI/1n1dRmb1KmxJfDO+vNsqrWmER39I
VzbF4PcmxCqNtdU/8xzhV7UZPwZNHSwt5oErk8W3N1iigB0bUkb50k6dNXDZWuUXrHXM/PcUqpsD
YpfeaOJJM8N/UOsKC73PPD7bcRE0cQ4GCv3BI/Czj225WfDfDU++tsXXlW7ZNNNc3wIiTM7XUa6f
EqE1AENX3ufVCRIWt9qeBddCTaac0JOxE8tX7TM5C4zrNXsjCC7JcyssgJhX90OnJ7O5IFFMDUyR
Of9Ltx4J4N3yPuPUp30pFXOsNjSI8AldIS0qBcR5Yn2ufVEKu65/M/83IJ5kFwoS1C4KiRRr7YYQ
7nhKDhkr700V7KRPMP1hTJtk9RF9KnFhLe1mzC+zyBjr1ZrmuBqUmOKmgyvjBq0Hw3W8lqTqzblG
uI7dNEpbEkqksm1Rg2lXQrJmXuuRCFr16W/v8GVDWgbowCEBPhYVCqKlzAhIRnw3+jNWSJZTxLMe
6YfW9nhZ/PDsfZQe6U1alwL/grZXItXfyL5wtwYS/DeAErCPuLNl9dcW9M1rG8uQOc/xPm6vTc2T
f5Kx/mydMFhfFuQD1++ECzaedP5sIv0GvNBk0u7W6bU/niDEAqL8ZlCdunKOVSdOryuIxbj1KeaF
rD1Mc79YLmPxb7gsz0ph1nQ9ScBQ9VIpCwm3+3pZfBuNHxC9+clTbwUy1DsqduhEEPUjpwmk39vj
TeIxPLAK2OIfbO3Z4i7tP0PzZfjL07sf+o61Ij1ykSQ/eUy34H/zZVOXMau0Q9bj4qKfQAcftjSV
Gvgrv8q0g/tmes5cba288f73V0N4c//EiaRqDM5s5mB1n+17rUdWUAksQ13Q2WMJ62hYhU2x4fkY
xggro0NkA6hs0QqXhj/V2iJVW3OP1cCAZ56z6KbRBZJpdXxukoV5O4CqD+ZZSiezrfTKpF7hWVPX
faIZeCNwDsUofjpr0Lg6DebiA2rGEi+llDY0MmZKyGDaBYEeCZ/WxEEQ0uN9y16h9ex3lRlIln5A
XIPUsoUUbB8OL9eB7//U723mi0QxwnhtlWk3VsX2wDgYmegf2kZRDgd2mu+XkEar7XwhmwovY2UN
EB+PDSwWCisJK22b7bzXwcVvlkFwVabz7PRC7B7YPvJTDmc2TNPi9ylO05b6wBHjH8sYenEeeVVh
FUvaaXU1Xdl725lgdOResh2smOQ9dUnZzPaGO3+yH1MiiOLH4ulqeWuhxjl18xXwS7U6CC4BGOab
vT2sAPExhLexY1NcpF88YakGT1sA6yPDKaV7W+1mJMMW/lUrO6b0Zwo3MvO83TuuBgbTSL5v1huR
cp5DQkmitjobU4uwcbc+idatSzgiMWFFARqDDejvWsORpbDzJlhCMEiO0JIrOA+LLtEU7Bb2gOm4
hmYmuZgYyFRvGpkrI0ymtL0VuNcnsR5oNLuJ1x+Wl9oro02cp8x4Xsn6xNK2E5xgL4pZ7pfc8bfv
wdzjbf8jwhLCTZni1oXusYSCxdp4syaJapeu5Z4va+8I58H4/VlwhOWfpRH73IB15MkrAz4Su/1L
s+trMKxbgHi/fBU3VFxEUbrMuT/hHvGFbdZfJVlo645AHaLYh10SPT1gRytxez2e+Sf0D+HZOkbU
DuxgmV07vt53G+oBkJoLXadfwpw+xT1LgP4POu3P/koOvhVDR6k1OgmZKAYRucySaB6z6HKwudbT
cCVICJw6I3oAcKiX7S6x2RvJdoM9GqZsxv9xAyu/8WAliNS+jsEjlRSiMeaoOjhztw0qwfav0l9e
r1v69WrN1wj9qKbygi0QjCDLJ3qvHJBHBMbpFCzLr8rgEXaA3t4f69ECEE8JaWD30M0jkgJzyP9d
I1N5r5TEItVPsNyNCeLuaQrEQgNQHZHwZYIIXLgvbdwYbya9If0Sbu0eOczDf/fH8nPvzS/m7jWI
se9Y0Tzoa6WqbERkmGE63qLXqaspJF0wmjp+CWqJuOeGJqwbfe0zypYvdPbA3pGCjBUt+v21z7hx
m1LLOCU9UqBsA9PiJOcN2oY47xDZlUFIbfZogun77atbRqbHh6S3NSk51Xwff8myZDpQV/XlE9v/
gd8flfnTMXq2YkVuAOTvvdrfR3USQ6A0nFtOdtVK6B+/9GSEZ/MismBrx3dhTays0zYycpFmHzyr
Ad4QzUwQKftvIIy6uRE/5bddEEE7YyChvP5T8M3AimJAKaGjXvydsCta3xogd8/Ngqluu99MEDoZ
OQHOIuvCuQQXtIEDX3fLvO/tHJnVzbHJ4bmQeD9+XIIXDKXWj5egzka7taEIgWrQIp0ZepY4950Z
JuEiRN8ryzDMPkFfTjX7KQQRrEc87TyOgZ2FKwnyPUd9ZLaEirbEL2PVLthCX5Prr0EPJ5zpg6CA
dIKWgBOluNLpHXLCJqN51IGffsS+0sgOnsVkhmXpJMzeQUxysm2HWJX9Tp9SHUgB9U+XgcrvieXZ
Tcf9AXfS/+82q34l58OESVNcdw4G8z5GsbONIF36vSAnLQtn8/bnklsVEl8WzvqecnZZoE11hiHZ
8UO15gY8D2X48OZ5+0GQFUnJA8qFuor2YiLTaYlpkLrUggk1yDa03Byx6aHmxUtqDmmPWJdjtbMN
a7jxNEmHR0qSURf8Q0D1m3wcnMfm8ZrQhm7iOQqf1P5yMN65nIqbEj/AvuLef5/J2RJ//+5Hj1OG
BqH4TwQ87RghT8who3B0pmQqnHPAhsYzAOrZy0sSnTjNRX7BTkhc6OD33Nj1KFHtIUryY0UQ7lyi
2Z8UsnBM/1s9gFmeD97Uzsizb1BumPz1mJqjXLoskYsWO+H8/qmCPNY6eCh8EcHShH71YYAMJ0bu
q+bfjr08o0iitTaJTMrs8dItO8xoHH5L/cUAKfiouKddbaNRc0GbLRzBDNf9FMECZEeOysjMOKkF
kF9xkX46SJlWnf6zfVP6HZ4vwHAPfUsHjqvbPPbyJfqUUZtg0LHHHKV0+FUspwY7hqy+6SoGO5fA
HrAneKQ/RW+pOH9ErWjHCAcYDBFpvPq2STWByFHpst9dTDA86FC6m8hUgrrQLs6rLq3l31mEygZ2
QYP6GETLM8b9Vz788qlfNMbwRSOlXzrrahnyimvIyjJXJJlamEiYB4wWc/x4dEhz7uhsMXDq1HWT
Pbx8cZAoWjsUqFvOfIMVdAuzDRgCL/CN5FJzaYSIr3iBm2nhJlt64KGr1tPuKuLKmPgbhbFEULkt
wu0uYoys7v+H4tSBp+AsrLCpaayvrf7ebZySNkb8iufw9DrhsEeeVqLx8O/ObrjWzVaz0lxEE5nb
V03H20aoV+/duA6omwsaqcVEAGBmAaax8pqXLzkBy3f14c5Zhm+az+JWvF9EKutww5lT2OJSKuyG
gCjuSuVaXJVId9IWdJGGMfuRiZWOJgGwY3mPX41oVQrqOuzivt13GrSoe7rxocr3iM5ITEPgJMZB
slR7A10z/i/PSRwzRcl6GHiLkF0nw+fEh/4bd4t7sT2vU4WAAzDt2yvxNbzptp7ImvpEauHlyJ7O
OfpbtYHr6g9z2NEfup2W5La76axqcq4gmDP7PRbKIfUZE/pp4H3VXBxJbTez7QBN1olCO4NXqKC/
jghSjV7Ck/zBND9jvNeJNpw/rpMUSzVmwA6ewAQUHPBvOEhZaEz8SFs9knEgYKabxoKBsJ/jKT1N
2NRC96EV+3nyFksTH0iKxWdLwNyplnNqCBdSy4UZ3u99abGqLj0Hsfs8ZDgKa19fdvgPy7MBOGy1
hhbwK3CN3/OqRJ1YeouziIcQ2Rlay7A/5/z3guIuLy7kIGwvWsK+2a2fgVN/AXzteRYbEkNm55Jp
vcU5FPXNNIdxwITb59tlrpSvcFXRZrPZxHYWJoxln780sGeHa0C2WvZlV2PhTVzYIBt32cr+JDV4
BV69sKrX/vCrUsHpm3VVpquj9+HLcMCtQvyAaJ6UIEUmSFp+Jc2v4bqmoDP2dFNhj+e97OVNL5Px
/YUUStbCO+voPnN5YC1XNXeV/gvYpl2UozjVxxjxP1ddj8xgkOzjbeihXJyc3hmR8+I+MV8GkguN
kEXnAv/VcVCXhcXG+rCqw/lCdoq7rkF5D06211AXIfwCYtQ7aEuE6X6SaVMdpKdTnTRGCBw0P2XJ
Id9RYAemX65V79ed8ZmJ1K9Tj3SzrMH74DCy7JAaaIU0yt+0PZGa5vIWC+pUNstKwYyLQStRAywj
h5eSlpTjsP6Q83xx+nNpmXN8qZ32aaxP657BPvKMhKzVobZyZZvk2hREx62y2uAlOz+0DAfOL5EI
7KL1iUuvy2m2wpeApJ26shLijFPJ2sC45ituhNYbCmJOVfKK+ULkoB5I9ogQ4zOh2Ha6z4urD4aG
2i7vw8aIXijWsz1G/P+8LDoVZN1e//FzeutzPnQyHUiHMVYme5DDvp2xSC7uVMnLbT2rl+VoQaVm
rJ8QH1J3x5XiTkxsCAaAvtgQoQIuRP0/7HT5v10+EPJLtOJHerP9g7xrlGRvWk6DVIbMiFfQZWN4
ygQXsMOb/z0XumU4JJyf/DeVF4CRYHNHCkD6lVOzsqIsODsbC2I1IjkLwI2Z5clzmfjoh9xSLwD+
RLqrmdQ1jy5xz53GaK89tEYffaHbaMWjtFFs7pKpuILzR1CYPhWw+FZqiz+fc1o0X3SVKMasb2tW
5YgAm/TkC7cXrzMfILtQomUJu+/7Hf79e/eWVFCi4xdZb/Gubgr+sO2cZo7Ct+tiVHCc5PdTbgGa
XmloI/X8f/oTFoj0N1C0/Q/vo4JAjqJqWcbH9Kuoig28IB2LHJuklWLhDd7MC1jMkHz27pgUIJ5R
atpM0rnUatvKGHLY/3Qvri59X/G6kYAvtw0FNH/pdHbzpEREbBQnJjBZbHmwsNCpAeakT1HP54IL
Lw53Fl19IJLYqWt2tm0a2R4UyMzbu/ZI5MXhnhJ00RNGoyUuETjhhn+jQEniS63ZnQ0cdlzhYm2Y
ApHcXs4KRGBmQ89QKxj7eM1hal/eM8N6f6rgf3EBTfslIFRTPjatZTk6k7AsjjDIx5gTLcrYOTNp
0JWg2ZpYVnotSw9h69mNId35P2ucO3b/ieo0FunF7o7FNH4WnV84gPUPUqbFO79cTL1dqWEyZvre
WCtp9A/VuGgdj6kEJIlS67/jh5Zn6XPYSALrDapIsHvvgKWKDaSrG6S+BzPlktvZJNPaCUST6Phw
eML/Gracl9JLGWpX+J0xl1RRL9SHB5tB3jHvb1AEhWR+9tx8XphgbNJe7B2PNZgbLwF8MRtnJKKy
w3HGLSJGHVjkmSla++6vqqEkxgAgoiVENaRjUA8LaSenKmeM6go85BGD76TVIqDuruZ6ITPxqQ8+
cbe/0njFaIBMY1rDERnoNENU3aQhZeRPez5lZQ980rm6iV94ps5Q9ypvtW5xTN+LpBgaBsy/1gpU
fzmAvUsgVCeywOcm6jxXk7e102KJVhqUpFZXqU2D4qIr4/fJi+hwvQ+frrQqU4CvvKKdtXd+gXUb
N9OP05AgdOuV05JiFG9w/kXgCSRmgV7IpogTB3F3nlMCEbVHtS1JZycPonXg0OdooZ4INsxw/vJA
iCt/D+kCxPUfK/V5eV7agYLdkbK+6gELcl3qlHTTnqy9GKZ3/dkWT23rawEXeRYOtJRLyzKYtJVQ
bkeg22UiZ/Oo3M0yUYJCA54qz5bq1P52fxZFNtj47482m82eBFbjudiB5wCcKJVO2FIJzq74P46F
QYMcJ5H1t+pRC2vweu2Vz4+GU9BALUgj0HLfYs6MtGA1O71TSsCWcUEeg+3HL5N8gfmyzi3/tsXI
7fqfw87ierXfXaqVhd1SN/U0l0EJaK4EA9JsDxHWpGQ7wSeEqjLfyhY3zFFjEUiLRYZdhhlcImD+
XWgBE3hJEmYRuaFV9aYe3Z8xW/J55yiXkq39JxbIKEqg8x7u65Q+vc/vaminMJYS772EdZMf0K2h
7on9dDnzMTxE9kD6LmLzsMi2bSoRwR9QAHMVIKVcHHgl+uS8OL5BNAhRzUWSmQ3e16iz2jZt7LPX
42l2RbN20ouLKVligKs6zjuwcjH1xjsgerQuuVf3ajf4SjOCIVRLBri35Qk7hjh3Ytq4U9vIYLhm
KSYEL8kEndAbeVgCWR4chdI/pL/knKbyyvvIwFoGLBZtT3gHIb/Dgu87dr8OiPvTm97mT8EaZN7o
yDL5Z36g/YuBHDXBU18bEuvYocNH3vTKXJV1OrFjWI+cW911goXZxKOAL0uZEW2h4Bhwl6d9Ep79
IdaENpfyQlX//rMawJFOfCVoFPCFPuLnM+h1RcmrKe3yl0VY/9f8leVhY/bNCXKTbilUwbN6lJma
ZZJ5YzUabYDKqEGoPBzQ6hq/HOk0rXuXh30C9WxBx8fxCbHd7TrZDL+17aQJNJ7XQ/nwgXj+BLXI
bHKO/QkBdxhdmiGn8dYPBwXKtuFYlFZB+pTa6pdktxLImAQGNKpx0zKnEFmPY7z4vA5dL1NBML5n
sAkR/yn9ce1DapXWnHSofy82o3cbRCwEwsCP5SXrvaypKZc4B8jd49tzb1nqvC2DKLkZBm+sw5yQ
V8A59ZGjAlNIs0NaFWMYrybES5pyfTi1WdmJYuYAABXobwZMIgyAvLJr2bDHxe/EjlH7VrrcSRM4
9g76jbcwRsKwt06rUIUMY3LS8rjaiGn2SmS9P1k47kgyEnYqfE4V2sTphGtW6Xy3Jl2a9u+2cI/5
SBcyOEqICmE63TY1m6lWWEyRorfEtkotQlo9DHso13Zx9f2jJWaJsTJguskV+3g33DU+4ZSm+8Nk
6zp8mQ/ev4B38KvKK9wEshwYfTPAzqjgPXjYG6nstMLyS8t7bMUtZ2QhY3FTLg2AgOuNcD9bVC3+
uPSNfJU1HjCtxXL+ezKRIrIlkHH2xpYrbxxODPg6jpM6cae7etqN3Og22ZxGwTRmRubPCQJfrd7O
Is6+Y78m0Wn4WLxKDAbFOuAY44XkUPMVe/u60Rla28TeYmNpHTI4bO/T9dDFtHKdE7AY83aGfv6U
5zkTRssJj3XI9fd/F+IjT6aai9IW0AcDn9/i9rO6FOjkmeRFK/5pY01LxhE08JytkK3J+pDzfOKF
XpImt5h2eiIRz1JXG+pTdkehWpENMY2ZY8ybt/znu5l4tmlr/9UXE1D7ewidIXvVMsOh9fyRtcCp
skcBD+w/HZroTPsLfs+g1trKr3zRdIy5E7MLB21r9350P/mrXj5O1sAjQnF1ZC3/tZv5bC+Sv5oZ
HPbSB6EMKlgMTJaCeZGPdcC+BXlNaMbxUlyUzgOTI9F9oxgFiIVDrKM8//DDjLPfLay7Sm5/YNoT
ULI5rMw0r4borF7lOXhwFPF0PqpFGzaNfdZjpHC19O8rkRzxY0k4G6Qmb3U1gaja/ZZTIE2OA1iD
+1NmVSbChwDyshkXyvEDRVFiOmWskx5RBP3OfMuYDLdDiUgHDHveIrulZOf2EhvwoacfMzTNChMW
3vrApZ6GEFUmCzN9IcA20QMNnCrcikD5X6bws5sQqMaCCpLYEaRDkWEvGUPFkCpI8NJDZbFpwsCX
mfMK4syTi9Uq9DHeDsF255aLwDNSD62H4CiVVeCH4Yww1rqSC6uxw11lj2WCLSWn/Z6iaOH6IsY1
o5sDDKbhBTofMpwsgc4RewlgqG1JDL325T1OXaotdrnBMhaziVEZIOlqPuaGA4H7S8cVMHGDFEEW
/5Kti7c96+ZfLSvJro/YLPlNQrWjN1zYceq/ltZzJfEdF5B3Kzdbulo1OtCFNGxoAsoPfo5kCFHd
m+ksLvr0kDr3zezl5BxqUOAfOXZe1LcnCf0Hh2dNVbEe3iSllyz7WuaOvURydfEb1GKtSNY9lQ39
XBIdynMdDs8cyde89uYjp+CjupGZzecranjIENXiitVu99kBcduGQJ+dSneDsDd8l6iV/YWoCVJX
6J3HTEFjX3bvNiNFWbIiQu4d7acO5O+Pfn3nkOwmvH/aRsKFD7NtPsYMNraCcGTxgfg4gzV3e0vv
VALZHCKY8wsYne4bFaQOPiFn+9rCzb77T6Y5zamBXpieWjBKoeBkOx07gabVgffdfRbKaGPOkrOi
DlcyTgBUCQ//7azZz46Peb48bAC3kY5iBnqk1YaLkxEjUeXBqI8GjpDs+jD+pBDI1+yNMFd6F4a2
M/sXpD+TaDjsKGO56+se/H3FmTvyygj9CEEMfX5AsOlVBsA5iiLbHBfw5pH0G3BX5qYGKZCV7XY5
2rJa+NSYmACGgmVBmD6RX8DEO9be6BWjji+VAljYkpipyik5mCS0YRiBWCkXKYjCzkCntsrwLBh5
P6sgG8lbBP+FWd63DHUBr9pABarOEzpXh9hHScJUHJcooX86GDUdZKMlsF7ye3dRMUzT1MihsPPJ
XPF8xFUwhyU0vTbETEScGLF8n+uhlatcn4dXARhOS+ZOqK/kpGgSlRnpHfocwhHFfVKinfENC3aj
fSYaOcwFEYDRumy5wOQP7wrJbtPYgq3o+IBeTuFqPf3FMI2jeKsfG07JVG7DnPnBjnMbq4yze+m8
0S36nXlNRU0DRaxSDeXP3SDTOE45o5L2DB3k2urI1JTrydmGhmNjPTn3mjOME8lq2FltmcgjrvIr
fekgVK/+aMN3vNKq/vS0nQWDhjeprM+FXHM9hWcYpf1oD3HBLGf++h9zIXFC6fIy/FokPasfZ53f
pC+USy5ldhyc+Ygyds5Ye0NBKPftxAecuZEZ47P6TKAtvyJ11SmetjzLJP514nQr2aw/UrtyMmVI
HW7o7C9LRvgwB3VUwzuG2rSFX3lR4NPEBVKQ2RLVA8F1vzzVJoFH7G+Zu+XztCfoiFFS5tDjp3R8
RSRlgqUAdctkXTwzQFcvs4FEyWeWm+zOxJjuNkIxaj7sUIlg7XW0xTTG0NDuQ1q4v7jKUc1p/FvK
m4jES5OJaY8o80HTESA54mrrMBbGtuN+VUKu9Sp+h8qp7q94fDdPZbNJWRPYgVzvJ/WLD2M+5zDU
PAaKrh4rpV5Ddymj92KRTrzzXA/+Sc+BplJAQzsvYS1i9qfqxyo1d8TTnpvlYjtdtBOzs9+96cB2
70i2tnutdJke+Dkp7bJixX+sw6hJ920RHjAfrl3FknKgydn1lV+00rXsyxzwGlR20UTjU18Q4Y9n
TCW7B0TdQyXBN4US7XatRmRVm/VfV+b18F/2RRNSh4JgRY/f7iQo97agPku7sC5A4bC6pwBNgfKq
wHw8sQJppQvtPGTk5jl4s0NSUlTQd1MQxt6aYp8GHvljecQw0CTRhzjlk7+9uz5QYHzxONl1GfBT
65Z1+ByabkpleOnT3py5ZPXU4ZUfe7vtyF8ZlGF+WS3jzAESpBHI7sqVy7r3qbbumIAY9VsN8SU9
UQjtGCUarFnp2k0xeN2259LHP6f7FLxlV73cscahnNqLCevHA8nC2GzYMGcZP24GN71EUlKZUYXs
Rd714YuxYP6LclHcaubyFzjYBkgMfIO0YB12w0vgUobHDF9QUUvFdizpeCzkkkv+0pzp3WCbUoFa
pOiwPhQgJuRd+rdxCjeY98KT3PlOPGe7MjUc200fXrYFKfwwOyU9Y5Rpy4xEhVflwW3/ui6UnMpQ
tuSSPhrmRf35ig3U27mCLAEoWPHFCJV6sSzsELyvGMulUKeizV86Ov/M8CagqmbmW0ZkxABcewOm
zPV/8L1sYwjgd7LzPdWVVZ+5QgrjAP20A2oNRzYx1a9ThUEqc5VhXDl6TviScscO+LgKcK1W3Pme
vhxRmCf+AsXTRMDyzFaEfHFeHzIjpUWEZTfbjqMqdsc7TiJd/y9K48eLkyhh9FFfHR/sP2cmxY0m
6UqyFJLrRupdZL1HVx7XG3bJlZUA7GruepDVfFX0rtQYTzyM1oRMRHg4kSG1iUp17sdwHE0TzjT4
20LODU8LvWMfwTJlH6mi1OAR4dey6Ju94+T4i05Gs8hV1dwQuBldfv+Nlo05MkT2FWBQjxrJbthg
acpDhJ6Q3OFncWTMyRGEsW3H+iiJuQYyFkIYiPNAOTbyOf+JhH0Fh0yIm0LKobrU06TQDVG7DNRG
LuCEUPTv8bzaGBOC2w8cZdcYOUupGitr+D4J8ltFv3GuTiZNfxYV1D7Oup8HrnJ4AS27uqoliNUp
yEEqoSDKAKZ7W5JZTAnXMIDIXfHvJAtNl5+powUDXHvn6K0R0Tno1hcJ0oq92qQyjkFgnLHNPMNG
ysrOmWSiM8Z3guN5f1y4TjeaVz/gbOSOulsKeW5rTyebOkExXBEKseAVBWW59Uh9pbbW5CIJhgyk
XZtRczdvditJ+GJ31pEQjxWhqDfyeH/vKXkPNRone/gROM1cwj/CPsHd4IRZ+hKv+Ma0Hu1eXIeK
iTeNpYiDAvM/hXBhWVk7S5ZPaFf/IZlBmxe3Yo3I/iCUmsn8TxFkwvnxzi4aZS+2C8cXWlJRrV43
3IHvsq8ePPFSp5ne4k94zQqGTIt0hmcGEmx2Vmfcfq8KSAf6ag0NUXrVw/I/++as1MOCurWBUwxR
blbvQs7IGSlI/52OT44YKvdMpSa0Tc1UcexSb5LLgSRyM9QpilltoDXJsqb3uQlFl52Eu1/6Plkr
QkPp40qG84YqnLn192VibmBJ/sD0zf+fZZE2iAktc7pk+kiycIrU26bqmk7KUKjZPNw1CG+AAAXn
ERt63ns8jlNanl3GGR41iniBcadAyQE0TjK3ezUNQCevPHpdKWekWaSqnEU+auSmmUc3hG6YdWH7
R3sbLV9oJZ7pfhGRe3uUZ1H0T0v36GSn2zWaf3XgbAJJNEV+4uMNonO1RX1NYTOY5am+DyQNLX/d
yxklKZcFuRiLukRS1mFdZHgyQXAIlLjaYaqDqd2V4F6QUXZeQe5v7SnFpU0Z8zk6OEARp2QH29O7
xEhSGHhrkMehBtJSFa8EFwglFsOe/LOHfXP8Ao/GuYTsmL6E7iDHJox85X9MbRSldpKjs19bxgQZ
9pWx5DMYWsu3xmOKUi3wTR94TC2A2vbjOU1AZlWmCY14Vh0XTdCAG18HdTvWbh8sMWFoDLAEEp7n
Zj2CEZOXFUJpdwaigaJu65ZdJq1Nwe/0Loigd+lmeDZQsfik6VUTUuJtdS2P6C1JjSWRi2Qlhqs/
PIPexMGMsPMHK8mPQFz5owl8NbmgrRUQHG3yx8aNPBaO63dVCqtdgIkBoSGoZ0WXUBpryGgq8ciK
cGmWY7NUSu9sJePffBoSFmQX+CbQIRrbRG433nWJJ53gakrHNIIgO0gMySot7uSQJXhI7l77BkIE
LKE6Cp3N2jeY0VVR9cbQuTfyVJlM0sQQh4vQHAwQV3c2GesPxWNElBfGY10uxkjXd5jrAWXEV8Oz
wkHDDJHGH+fHu2TK9bLxF2hieD3yt/y7j6fl2TZ/yD8XWscwOy63/yR8A2w+oy5Xs9iLJ9OcLsOu
8u791aL9CQpOjMsiNZjWL4WNXpp9tb+EtraNmUUNyvI2WmlNm28v+fkFGibN8GEe5pDhzbgQ4YS2
aOtfsgHxY+gx0sB/aXCvQljDXG5Po5Nd72ST6bm1DjFsIweX976VQtBLebXMWgwf6NltMjcL8Jw+
TFL1a9niMJ66aCEjwN/Ss3B+6P/+YNXRLiS4iEpfHPvlDhOwuUBENKygCnsgn0LkAYz3lYRckNEu
qE22K5T0zxuOu51H2zZsAy+q/wY/joGi5pQWED3HZtRQr1r9fESjkLb3hbmsngHYlGYDsJCJS+dn
ciJeSSdo0YFuRJTxk3dG7KSzcmZ44fKVAfNTKoZm6MveZ0THN4VgIZVSk/OCLNCACZ0NTs5IRWEY
+yFV7RGa+60PnA59nmtRQaT2BzpK2fMO0XW75oAraL5HvAP7kEajs/YxdkCZKmmfii9Qw6D75mw0
l25DrviNdFtNyuqoGZ44rrud3PvEAxdj1FKb2OSmuy5NSkLOThKGi94fABKVQgeogrRB3c4kUUTf
AJcV6T3SonnI+j3I+mrFNe8P0tLZ0ywP474pe6360Tp9hcg0Sp4ebmaE/1lhBwhpCGLv9V8s5MqV
/r8V/TzMvy7Z+2e822o3HT/rNkH/u1sGaxabkMFu0tSLb7xYhKBXubKoN/TkmdnY0+4dIvjkChKc
m9xjh34ztyZjB7kEGy9/Q1dtWV8HWkSMBiacSm6fMQ27pCldASW1N9k5rdozg4WI/maHMgeQzHBu
ORAkIPAaleONUdGSRMaaXqrEnyM9E8oKAq9QwI344w/UGy1IZPS6nBQh1kzTRLG2npDUBhMay9ES
UDRWWdZI8Y8m3Q7e/1zJjz13Ot+ESUJDrIKwzxXurBnw80IztnW0+0DD+l7QsGPPk5RYLYLZH8TY
nws1lz3y8OEzltGlCZaIGBsoYma+I+WIQ2og5LRwcjORlq78ids0BXulzz8LLHw/RfuLJSm5X0wB
UODG10X6kev/nJTHcBjXc+ZslO8MQtB2TSyC9m+dvMbfVDywfie2iW8663XUXFnh+LpT8nme/7M/
2uoHoWRkWpxlNtgOdtaW5qNLOfZcUgoiJZyQMi01vUS9DJds/8nYeIRY8D8BXAdf7pN5WaAMgsHc
74ZHSIe3nMBRfUZdo3uq6gm6AO304hLuX0WBItkGIPRQD9Ch4695Ys+CH90DGK8DmacetX0ccmZP
qXj7ehGjl9FCAOUhnkMVl04vErHRRUS1SCOximHQRmGNNMaGTc2bMMa2DqJLk06s4pGCnKzXGpCv
w5zvMhyDp+V/0c4iJBkRJ5AM1TxLpqOCahgMzIYg7OmWqJKN3nTbWFvHWR9a+OWtvNu1ZazQhlkN
NqE/5r9Ty0L98KfQ9Vyd314DNUCIYg9UhyfsZfz7kbMefxL6wcvwYIWkdJ9ztCILWz8NiWbOVgPl
18CsZV02MT/vGoUcP9xA+iqBFKoolQbuG2ugtk56by4fpqVaixkzVy7scvgdurrbVoH4PlILYY2n
2uqsD7HUmCvbVQaIe6gt+OAvlQQrIqT8gBfylcekmE9nvxy4UkLP4eugBCUIiWQMMwkvPQdvh1Db
ha+BsuqxtRJ//o9vJh1xng58DkDSrRASfhAEtvSTWXkwKhR0A0W3GieyMeZKmhghlm/S4jiOWyTQ
+9AvX8aWpGu5l8hhXuxd4OFKnVH3XlDNd0KD61GHeSHamcw7kEUWB/FpbhImg9SBadKUug+hXBFM
wCKmHKSjybO7//1NQkiy2/mMQubot6w98UE4uURzDyJJp9E1ec4p6nMPgeuJ/iAcOFfMnMDJ6/O4
/ZLG9YNMoTWH+jK76L/BixirmmfKHTLM2FkcvWUaI6muTiiLcY3p0/0w9Qaph8sML+7yOvzNoEDF
+whbqRCdObWDKa9opZtqqCMAxa4/ySfgt6TdV0p3OUs+8o0nfUydCrX8arg+jip8eIDUkDipsKBi
q7+g2WopnGkjMKVVadOM1qKEDUd5gEXqUbt3deltmnpi/p0ZtkGcgg60GADjsbpygtVhDGEvUrlY
rskSD9J9Tv4t+FOuyc09MwrtCvEldzpC/eW1wy7wzHTnbWIKOA1Yrh88IyUjmWQAVRrPNvw1W+n7
bnZc6PuJIDi2mYcnerVM5h6wmSJBIrzpmq0hC52XWofeOytLGoEpoM/qWJ9y1KpZqgyRl8aF70O3
lfoGiaT1L8HygXwHmXlOulivJ83s6R8WJYzYIyyl66PqcJ+zkeGuCI8wPPJsoAuGvCH2oMmfv3Fm
uoe0k1yshLCiUHLjRMrFULLeK77PX65wotifoyJDQ5cZQHv4rSk5YugFhaoP605sAMKOUlnqf0oW
kd+xXgrlZovwi/fR5uTZFesjg1a7LPrXr483UlQYxpUfOcC+/ZII8xj9hQqyqGigrvsMS6mxDU5t
us2awxkvxiCb8ujwVKFNVYmxS7sOOkij/QC+cTPbQs8Q1sG39/fYWieZAJuJF4a0CK6EVnqhdwRg
45tFuCzJyL9L1dTJ4B+X/ib/M8TDnMq8QcEr/LUHG85L8t05ikqeeAxC6hFoUhsUAxajuDRLucNe
1U38NZqMHiT+S/9ieFykxGs5jiMi4HiZZyGww1Jhfu6GKrqo8XgOhPpf19yZOhEQlFkFXscYD5f2
e+IK+rohh+u0BJHLbmDSiJj8yNtczv2vlaa7nsCwY3D7jUQfREQ966jKyPmkVo53F6vKVSdzteH2
AkN/c6jMwwMzLHmsGu3+CPh1IuTH8x/udNen26EdxzrWJASVJAwqB/SgGsxHMAnEk0Ew05QV6eyx
dFd2Spi05a43W0Pn8Y/Ksz4surQnZAaZhBjBMUgHdGl8kztO2k/geDWDHIyJaxOkAF0IwZcMtYjl
pKccf5U7PzUIHTUY6zYDxhKC4NzP+WPHB6R1c6e6nbJVKJglRNIdRhp8gEV3UD+Ya4TU3PygS4ND
/7rjFWYKVsUu+HaZwxnNrM/7LnNTI3UIMnrCLI51HBPl+Ccb3Sp5Ju8zqSD9uzEjnwL0oUuhzaLG
4prdcb2XuXY2KWQaIBIxTAQtNXlv2lZlByxdLnDjpGyFL3mb13dlG6fNAc1TsD4IaDWvrnf4VYv/
FjRkM7pG48xyhpxIshy34n9nsmTHYk/nloUMvUx52umVQtXoFxXudZmu9fn9iWA5+NiqJpgoDSML
+NENaYmVLFWu1uU1FXXrKBeYv94Ft+TzccYJdLa3Zy4WfIIELFwZ4w1x65CXU+WDJjETpxIwFJ8A
49VjE6cgtl4/TQns50b8cJHBQ0L5678vnlyfLlcBCrnRjN8dZzayFm8JX+kkVK1Ma8dEt+kh+qji
rI8ugdzRqdDen32bxfNZEHlllFkkOvH9vRDnqd4XbJ0kXUoLB++s1Ybf7/XUnmqpnMZetBwbTgpA
ELgWw4OG7bjJUn1yyUEgOqObUcEnZ84HxgYSMWtd7gSE1RhPSIlaRF1Xqb6aoE9ZRitx5ma2X5v7
pqrsf4fzQsyDuRv8wUpxVQPXqqQrFCTrPp1pltyhBoJgf0qoksv7q6hMynta+aZXS0rFLveq1d95
giwwUz14i8kYACmhCtIr9wndcpQP6///yGbmOWIvUBmNKNatNrQk5SGFqAIW7H34xfCwJF/Ykb89
XbAh/xjGfE9dyr1di/IlQjfTNAGpRelE7heahn538q7wXRn1UMCGJ2ffOyBs2IbPFWEqKWuxW7JR
bLUClyxsMzPB8lltkvv3ShU6DGToHpQ8BDMm9xeGSNaLl67nozoHs/wvntjsQpYVxiLpYbsSWZnd
kVn5RiYmpTVTMftnnrQ8qRT1Ip1OvU2p+11SMmUSQAVaNz0bZS5A6F4upBQyenlvWwfxGI54bOIA
EZrVwdBiXfFlQxgKLS2EGsYfxatUcARL41FDec9q2feHkVwctuTr+fQR/BO7vYDXGcc2tmZsCrnG
uAZzwGgXrdccpRYqVcc1EH3c8VefrXntdUKDt65Ul9ZQgLZAENf6LcfjLhAm9M4Quj+V3k1fSYzQ
vzYsNaIoYhEl6bf8TbLuPYuVnYFQ+4QZBhL0xpZyWy8JinU4ks1py4X7rHGzI2qkN6obf96ijZH9
hysbwAe1gglvgpJgqsQZ4kTgnL31tuTjH+d73bLTQrXV0k0fa2xXLMfCUG06Vd57RrMMsEBaa6ud
HNdj4jINfvGjG9P07Ce/GOJisrwH5SFAiJX+prXViyD0w/Jbn7CoG1PsEhagO0bc6vCJmP+gMn8D
1J9dXK56a38aKSfAqCjIcsOsaPlOsBix7OonZluG0/Yx3ePMrrjJ3Pm+83/km776MvwHYsQbV80D
ahuHs7XBF7PHmBXNcWI52tkRWHEQkC63wm/+NYEmOHPKen0UnAODPBDhn1SOFkLyTR9w+hJdI2Ja
efUD+dTN24jqN7HnrZ8ZAu2D3XZoRe5qdIaHWV9hoFhaKGjCLzgHJJJvsHSZyMbAgcVSQZuIyasW
2UStxsPYoUS70hG7xBVdDD5Wch2tKSXExPgzVa5lxSkGqqXAa25fByUioJjeJKQWeas7rS8wtxut
/EDAUW2MvupESF4v77M9ifWmmuMnvAeTmVWRWaARXjmMnpxAgSFYhDDO6QYpYcYOEVEM5FUG0qtN
LLAOAtIR9Y5IqqquYzTRqp3Ei/z8giAOC/SuCKZJNbm/iXsUbiZvvrepn3E47ETf2Fte8VnE6ctl
0E9pSXJLCeLNH8eh0o8x561oQvdOi6URK7DYCj1c/dEsksEU/NCenz4qfKEV+IgpyWTnCIdAOe+V
nXC3vrDew4Q+tsUVkFq0EmcGomYulfu1Ip0/0IilwODz14mFlJvY/ddd0LvoNDKPxKIOdOwAfeLv
AXvmGMJEzLcG2dmpy7KTt8XLNkVNj5mudCxAkhe65/SZCi9EphsFD3SFELd5L2D9wBpyg12PXl+6
nC8E3gImxtIhlU4J8R/YylV0S3xnRWNCcB0QQOdM0VAVw6TZ0YW0GkMQt6STpPFce3s+zgU6vDG6
TS7+MgfJhOLFTj/MycO+unM/mq36GIVYY3Jty4H4yVObk0aFXaFpbyeZZ5cBGAUrtyua7jbkJ1bu
X72W/9baxdG+YpY8WXyuQ7A6Ph/KhgSWVwlJRUHW26Ip5s/TYBRKhCycgN3MSxAUtvOX1dMJDq7S
4UeRzj97sfbWJ3jOOga4r9W6UWlk0WyPR/oSZh33AMPKqXzSi+6Of3y1qC+xS2kR2ZLkzg8al5jy
wLUt1h884YTFmoENLZLXPooGJIHy6/mkVfDFDIgAJP39eDIPjOr7kviPhn+C6NaZoqI6e7GLpSS4
RuUPTP9gXFELMnEWF2bmaJDpxz0PoZlcXjIjxCMtSA33CqF66uuZ2LPqfopNZgD5/Z4DKUkbEN3J
gQTyMHO8CzCuVbbKIuYi4shZxEUFNeKS2RYRHgBgikv6UdBxDPpnwnBB4eBskk8Hv0Qi3aK19GQ+
4B7+6xVp4RODwEFoEw44VS4C74ym1Oyt42SC8dNsdB9zkGJQQzdWXyqFIty8l4IBHL+ckVynBC/Y
BlibmhGzdIqXv0OrF3dQI8vR0UBBIoT0rFtWZH0/QmuWpzxN977iSq++iIhyoTEPDyS3T7M10BPh
JTYhDGo7q/K0fvNS4/nrMtFSO6+yP6SNOvkdohQmWSagWVRvU8gZsCD0t/Xqs/QqzO2/OLwIy/77
VtKw12b9V2BoBalH/mW4tQ1DfMrOx+JN1QD5Zz61pk3GUr+WIiEEyBRr3YmwaDrZBOELjj/NYviB
SYf6ZgiNIYPGCTnC/Q9983St4U+sxB9GH3vwXL8DBnKdadscQRDpPcaENHn0SL8hJqC+b/8HMnx9
LxHXxLasItDzzwdgVNmFqXox6eTzkneZ9bSd9m63AVY9xa6NSShJueSWWh9ruv5bA4v+yzQlX9EH
HYJA8k+4wsp2KWh20toRE78JScplF2sw1v4g54sH9zQ+Nu/lUnuTvdiRONix6ZyNp6dRzK/tuExk
iTmGYXDCdpteAUPbqGrnf5BVRsELwnsb/BS7o+9qJaymRAEg8Zuoo0g2+rYymP/18qJDEOTttcJ7
ZfOILz9LZFMyllvg5/1zp9zKcJ9uUkbbLIXIbv8cV1CPpcINSW5dBeu7ICH8+BN/60a9p2SlHG/o
uLWp4zT8BKlBBkyEp8bsQHPtjicgiVGurOFD29zLo7cWhR4731SbpapI9zzbug7qTAgE1px8JN2L
gtipUpcQ6WE/7fq9sJQnTOHoAfoJKezZ+RHA0GVC8wUZlN0mQojEyGXkLjrOsO+rcpwPcZFgCxj4
xyQjYApHKO1gjU5RaF7Ff3PucnZsMDljGMbyHudGYIRlz9FUlQ6YcsfI7kwP5eu1eCZOBgn0a9wj
db75TrfivSCrgdLceWqupMfIdMo8q6+oN+bvRIf59y83/bPA51OIKk9kcuu7s9KRsM6aiEv0UTtL
OXkuVsjUb48//mDAQJi27f092MbV4GwHW8kRnCcLOws8kGkKpZaJC6fvrAHoktYHzWHibQ5rpZWh
YqzF8za64UuOaCilybSX5rSgyAseOLvVSypTYRJ/5A8TV2HGe3DnVHVVy0RRcx3ZTQ/9RkxG6YWe
JO+ssjPEWL//tBZc9X6ZhujQLy71AMCO5xYHuYf8tymACvZzaiVkA4esi5Kr+NNzyd9QevuYsbQ1
ICCxs5/8V+E7qAJd8lufZGumykkNR0lLEy+JXm3qJ5/dLPnlv0GiAd5fBs4+Y9PHyq45B+sQrZtW
HJrypozyZL8ixRE7qkv7c8jj2lmJbIBHwu+N6HaMIBvbxE6qsnSIpecPZ3eN2KTvdW9vzv7rFm0z
S7ZY3mt1cjpE8/lWA2LdNa2MwRGMnaVBcOA5UKzJsUiYKNgpb+LyuoAHVnm/A2EEVsKTN0YCz8vU
nk4gDcXIXcsuxHMYb87yVTjasWYolQB47ZSVgDrw274blBLS7PLhnyriq+jNNy2Z5l2rDBODpRyi
OgXETUd0MieLeNH0rHsfVE0VBsVJD/s03NnwkDxgqDiOUF52xjETb9rm/i74GoDVIWCmpjmILwr7
Tldpk/ZQ+xSvnmx1T7bYRo4jJctQXwUtg+fE84ai6bQRi2tj/DhT5urMf+iigB9m1ZMmyZSoVLdY
LCFZvtX6VQ6Os0vtyuGOlH7+pjL5n83slJrUjw6M1fs6nVxvc0519R49iHp6t5MSYrzLcYA7NRkA
je8DKDpZTb/e2XrS10PpSIJxbIkSJXYwi/R1NA5R5lfjEJlzC4ups6dArvB8I8/zU7erHUDagNmb
SkVFsBfjMWuOTLH7NoLwkcS06lX6IdYEyZV41IELdGOqv9R9o68rfMEDQqWjMO1VRepRug85oyYD
h/Qxt5SdrnNlNbOmz0ApNaJZtvYBhAu52zTlz23hig3cOBenniuV1VHNtDKDI/3kBOpA2EckwOu/
ZzDwUAKEMhVAGEkOu2QFV5f3OmWRsUBl6HPjouhV8MCuyrLsiU1MrGEFjuWDyw6laixZpD5KwQSk
PnP2ETW3y3g4tgKsU8CSw5P7oNSBRc5KRKywGkBor5BBRCrTJDToBmfL0jfTAIFwr8vaMXYsHCU8
J83Xuvb2yfhE3k29ktA3XEsmYTRMzpa7VizoswGB+wvOTAaTsT3R/t0oFjkthFR9Yim/CAkpD12t
QIWF8VKL4raKn+XTDE8xpIt8c9XI6GsOSeIv8cGk71vHgdAqHB780M7bjfYERKFqYP0VHZ/H6GLL
TSLbH5+ceElc56lDg6tNMyUmpAMdHHdJsFCci6otjAEJHVd0nGII0WO6QwbHLg6DaPn56ovyW8Ca
zNSb5RJWZ90+dIvRNP3bmUHuiNFMT90yiyWw2qzITqa6mPFiOMPO8dsi+MZ7Gk/KVlmfbTRneNbz
GnoeqmI3l6cpLeOn5ExzNc5WeJRU4x09LGgpcH3yyG2OcIlMPIk+nfjm4qtTI33oQJh+NLzAySQo
QV9iBeb1mgNTtM7vy1J7osKWqfylg3zvkPnWBLLgBA3e/JeDtwlrceGM/KjdVGJ7CTJYme/JF9J8
kMNTqTZfQRI4Y1BWaOYd+oo2rutx8hbNV+p+MgJvvn7Uh/MNtyffvkWz4I3MxW2g1wjEVJXuo0Ur
wb5E2GiDIPNi0KIys6JM0sV04CrqoXSwmAOnP0EFpyWYfkNCvRtnZHb1VeYpA3xqou7UWIurt/Ew
KUkbDojnD7GjMDQfF6xIhpjgqmOU61ues69IvcfXiLpe1JyhEsZ3W0n5RRqKKRIQPhGra8l8aFut
JdR/94Qr+FQtiGe7S2H8NYGjjx3aNQY1qhyOA3oZLNS1504dzr3A5U3CScESOythudH0YS7gowRe
OZXghzZVyN3TixlnZGoLWhlo2zK8ATxltJEe3ntz90TTa6lEzx30+8AfzgjwT26mSR03l+b07GqH
weSzsb8Mg1idpBtuKyDWlAvtqRn2+Zjjl6UZbXSqj72kbuUcV1aIVQ0EvIJmL1Xe+hQty4hY4ADE
sifl/8AWJW7UYDf0NLXq7KLufSlQ9b7Wh5uaPiyP2z1tYlI82zlNhJn2tAH0Q5hEnHx6MvcSYFdS
vBFlcs/7/ybLlwz/67FdX1ezFR9DgKBTuALnEDxtnvS0PEVoiKR5U7/TnRfj7rOGdsUBzO17eFOX
uggVPFFtf9+QkdefmBOCLKtwtBx2zTH4oDaqg4FVxlw7v9TnSdVgPC6TDxSoLpi53keW192ieEOO
WWcSPv+9wQq8PpNNBMuAljXS4VtAn0D7eliadgiymamhhFTOAVU860kkm6RrzB8rqRRGQQr47msf
qZcSxPsbBNvuEJJdQiyPuI2ATnRRt6Ofxl6nx/QwSBglKUx9NGeZs9zT/JWYUqKsxm0EeV8tfEiu
VMuGn2rbJWpRfLiV6eQSCDGQW2+GCW3E2C8qloatgynyPY8GS9ATRZgDHSDBcY9PLbG5xkkqfkUT
Z0j0gGq/juccTccyXNz3zvI7sW+I+giCt6GSh9p1UBkukf6A7KvASXGUBz6BbTz5wNIyeLoWUr+e
8xmmLdjp5RW4x/DinUBMHM0JjNUpLpDMPDRgn1vt3WCldSwa8pBNge6MlwU36BzC+GYkffdp+DJc
QJe9TXUGPz8MyKzmpZ+y1DD9/lPpzUzxg71hF35crod0a2TPWYeY6J28a5YnfI7Ki4H08QwWeh7O
5+JI68+j09aGSAi94izYN3qvc/2CVmc1IWvuAgpscck4j/3sE3mWlF3TTBJPwuAK/2aAz4Lf2HyL
E7ndFrlY8hohM3vKRodCPtHcObG9IuyoCq+82+j7jIfmDIAlJlI9u1IjPvgBdLoMUtw0whkDfs/Q
zCnrNyY7y0OfdDno5uNcV38+RTL/eBulMNGI6qKtc+Z95spGQr7ERZEdVquXHKw2w2biiOe4vb5F
Kbaz6pc96JXSS1lt54Z3QbRTQqLmvjzw/fG+WK6OxIsn2dKPjGofiafCD8SDPdGoWG7AgeWLojZV
2x/PdCDn1NRGIvt8FAOITU7Dea7brxoX7g5qNUEZe6cfhHl0C18s0yUmwRjGSulmirKzcqNYH7UB
4RReCT/rlzVo48AIxeCZYbI8XaL3kVVzD+O/PGVgxAcPpo2LrFgOTrvM8FJ9qdLwcsEFjMjqoc+V
K8KGa5+iRXxRf7tTzWbc1onOq24s4DhCpx72ZJTZXZIn/1bTC0yQe95mOD6ybycdsZpTQ5WKSR7M
gp730r0pXV96Mhq3cS9RBQKkUsoAyz9OSO4KYqgStMmuNN9QLgJLWK4ffU4mTKgnL/VCJfqiXhDs
5GN6dYMbPOKEk9Dxy2sPl1MQg/ivdp6AamaT/JWF3t1SiNQKx7C80xtcIFWzrZ7amT3XfN5WDx5f
xP/D+SL516sPwscpc91V+Mzx5gliA2MVrjIIoQ5ZArTnBsBS2JgxVRT5pMf3a67XyyhUJjstt0N+
owALVg7vjWiTgcZahdDKD1+gwV/5PIF1u3y1pcED9fFnGZAlfvRld+L9Arx7JIi5pu7/dts8qIuX
9xqy6q4i2HqNTuXr6FHMaU9eHafXnCLKW6jJtJ4CP6NNdS9m65UvtFObqOw1KojGIrdXO9jioCoU
QP1yLtHXwyIq8R7awUwZWHobhk6kPNIDE3IHO0hr1nMAHk6t4nHewEtDXB6ooVgB0D68ykan5NkS
BuEUrA7ssyn70Jm27BMJ3nUJTPsyqnwRxnZmxP+T/YWA7PsHtAdFGLa86dXwUTVgjFYCUS+2frdi
RYd360QjFqvuZvSyk1tdEBaKwFIlycilhgtIlqdqL/FH0C8zXJa/yBKvKZr/R8vmr0W1JeU2pan6
C3oZFdgGyDSmAWbQsriHg0EoKzJLBAHJlOlfAT2JMy5wrWVed5vWemxa0phRniOtWZW+q+s+5gAI
+FJfyytVIZ16yHXZmLvDPhFLlO2iBkVvyObsEXzH7u+YX/jMPm9dzisz9QkoqKNCIh4ZHgPBcx26
+v/OebdLvNBJh7197TH+xoLYdAeZAJ3uGVGSmXnFRrEKSh083ij05r2WUq5GjIt/0ml7VBGdIHJF
WptgUyEvReZhn5vA+tYn4bCMRRZhmXQOkg+5J+WIMrUbP9layEGe+gAxBBApqOopJv9BcORIOg3K
42Ku6RVRA4oTxMOeWB2VNQ9HUit7Xi9stnzVNj4rouR3lkownr4EgnqYCVb6WOYmml3+qelZESQs
s70fyAGlSbd5tTn3JC8ORp3IH4aRtfzjL5Rq/4XrGner6myAK9zZl+BItWMX5XzuOG/RQfzs6rI9
dSq5cdvr322h1da2CjPiVbwWAA8rNPgRRCx1xNDAehtTpjoxa0Ogw/tlpLoD2S1jgVlog2k8XI/3
Ms7eRDbAOy39xYqpZr5PbdNAF/4fJRGYbOE3ooWiO0g8Q3gvCuzfp0Yp9cCJp0hNn1WAIAMMfo+k
Gse0hX98hDfPiPBm2TkY6Fm0lcsIDbLeXBXu4GkdXepTzDVkmO8NjrjZHvFz8dhQzLcCytGRg1Qg
hzwa0wDHHRCAMyBC2cJuqFQvjv8NR5lvzPoMM9IfXWL3LV6tuuY2pjp0EE8s0oqvsEUmyJVuTIBt
zknUWoAvQ1/TK830HkSd5Wk0Nk980dS4Hyf9YlM7I9RFruTxpa0aA66f5rDvFm/SDrbFOxL5AXoL
FB75jU7w4vFdPJrBChA5lUe1FaWXKwWtF10Ab70O8Wvgxl9n1B9CEhi9b104hxCWVjSsgLzDb1Sn
f/XGfDtdYZ5How/0kcNkwS5lcE61tayGIuoG0wy3cefC9JMKYXh/69FYe2jYnaSuiTLfwp9uIqF9
NsYyBFUMRUFmcdAwLcQ5hLuBBqOS8kaGJOYbBcEzn/b5qEegBWHtlRkeCNKtEXxPbAjeVPBk8GGy
hlY9x45ddPkZdGTdrhEDAsGKh4XSNBzpQJ5qypOunZx6B48Nq+iAXVejHpik/g/ZAo8vZjaGsd6G
Z3pE5lziRZAs84XPkuY53vArPJIUyg+mNjwPX1YlO+tn6CLSjf4eU1nxRaE8KlMzoMvviuMOwR8z
fsX6lX9S8pebc5K+KOU6ALwg3RYDEIPdTsB/W+W8cjjtqIc6Ahl5dy7PSqUGHY+F9UwGXe3qYY2D
zzD29eX9OOe6cvYQYDTRvM3GUyJ4QQIIxKnDJCH6NLo/m2XUFRKIDkjWzC8mEBMrogMDRzl998QN
q8nwcROakGKqoH3YtYQndMpVmWGzX4V4a92zEUC8ax1E5eNN7C5VcyV8yL2vdlwhXwmoh3bppuWC
Gio/cAqmhtoJ1F7+aUGqiy7l6MRSPAEcgCxX+UfTpkBbpo4NivYw7VfBjLByzQfffgV3T3M8A7QD
hWi8hkOuZmvWpAXRZ/Fzq8MWqTy7OtsO0Cvxkua8MPNK3xoZoqQj/f9Yk2P1bITM1eOADcGM0Bwx
pTM82LiFM8MFqh9NBONSnngy7qGDxWzi5KM5w+PX3CdM/YUTbm5DSPaccNe1tldvNJqxDLMlqxSx
WB+/Ip0ioK2R5n2bRu8cJTDhsFgzTO1IvqTW8H3io3730EBmQh7LxlG7tytVildT/L7dGWPpOFWc
f4v1xhF0PWq7/1iSRKyR2R47NZTOgeWSnzY9GMf8fudLGX39Afm0nIas573Agqvel5Q3zqTiR2Fc
XKbp73sctl02Vf9feeHNqIN1OS5i0uHXrVYtLZ6TEeHNsEamsPbj0EnZtAxLEVQiy9h/KyE0Q9Op
HYla0YECT1DhW1CuX/XIRgJqEOmlCEsDC9rThbL4EhUaGgippBY3x7xZspuUObwbLWMzo+fy5Oux
11jnvcnwVkkU5HcH1LWAsBZlZeqMXtD01JQ6r9AEIf2GlotIsGxGB2uAkEf+wsXCSUYr177sZ1Lf
yBHW9W/SvtcTq9doFvFKRwe4v99+eaVxPPL0/Mrr2w3wh+1aqOVGKrXhNXiDuS7aMVo3/hgT8Ziu
bqkNp/6w7cpmi4j3PqLg5ShJ21ryOOZ+jUcbi0bZOtrRQy8sdDK7yyZeRly/tfs3aRputNlGZs6B
hTMsa7KaqjE3WyzUhQMhaYfqHOxCSy72j95iuTm+4HqDT47qxR0iMRkUL7H/MJDxWxZmDB6c1g98
BwQczE396KAD5WC/lL+tOMajmBHXvVXF6E8N+5vE75PbyGV2XAuf5GO7fFdbUh7YsTfyOJtOdPpC
lMHLANyt1BryV0KpG19xlcc1iSOFNGdbSwJtSHeCmoZ85OcUlyixJkWXDcNMsM81/4d3RP1eSQXB
yTMzWguRPBp7Xt3ms4gqcheKkKKddQc8I5OyHxoLB+ACFvDSYxunCM5uTZCKPxaRnNPFrBg28O2P
0QpSkzFgiUMegHcRP0V+h3rfr1mEfHcGZBJXXOtJJ0g3NIxkgEdTF3Z5oPN9fB1Pb51Gfrcvt0+I
dgr6RnhrBwsMzjvHuJ5OKBXL9qpcDi1NGJKmpG8bVC7FMap8M4BfRLd7kXy1LG3sKebR/FLcvnth
b5yB8W0H4msSUjyIEcnTNWVflwIVumLr2wU25pT5vRcCzzU0P10ODRyNB8+s9SOHZqs12fq72YnY
q3nj5xX1n4G9Z20KZvHGl4MzNHryPhLW7lO/8Dbe0NdVLY23NFktWKsNAEdzf22/AwVBxP+gEck8
vjw6YeeFj2zyRU9xDRYEvHaEiklAGElPKQA7rlaPy/cXOJopHFUs9lhwsWtDqMEqFg3CsxnyhRRn
mRJu7X3B9d6EnYin6TIzsnZaHMc7wOomaRs23dMI5LIXyfiI7Hi4SYM3c5R2WkDJoL4v7Orvyq/e
J40BtU0rD3N1Ixh8p7KaK330lu84PyaWZVxTcVjKM6PBvD4hhL0wNwxWxExASly9ctwE70Kntdym
bx+c1WmUIM5KhDl5TKUo6FPR8V0zztEfP1oSvhuxEGWXZi3IIUTf3WMA58zYGLbe7AHAYKyNAeKH
XnMSFqIGiaZ2Xdw31QqGJRDS8h9ltEZLg6uxLs2u+OSUw3dRiwMtBLtXZMpaUbKGAgSiEbQJFyws
te+dm+9PdeP4rTIJJAEJEhivgypJUMwqdUVPXlNlVkcD3aMcVm0FsgY6wZdRHAHC5G0/sRWQuxLF
IsKhoD67bAlVM1Yo87Z/kwB1qTWRiGf23Ox6Ipp1X4CC8CyamL0SqJubN7dacI/LFbReyC/8Xhzm
XIj//n7FwWIVnemtDMM2WXbD9ssYIdRO4Ze+zpUSIVHJhdXfEKOk4wevTW9FS0Nw6re6LUAND580
9FR9CVgpPO2aa4CDNa6f1QsNLSn3zMiYeGauExaCeobPeP1yJ0T1Pl0Q6dPSk4gGedRq7xof/8Ln
KExOaLjukZQSXkqtjbjHRHdbdBLpamhtoIwiHS193B6G0p45mOLIPD7CKw081DTEJc/Xcbav6pf7
tiS9tujLv9DWhahAdkyaEN796jArPiiGmqhEB/id59bBVZXCxccm3GAS6TLYzlmvo8iRnQNRR/Fg
/NSRV8NirpVl8lkwEKerVtl95WyUqLBUSjfIdTBEpyC+/arzzwR5HAaN9BUKFV3a/2KIavzLt/GZ
op0JHGvcX137li+zUhvq+cNyCrZgTlmHkmhjzqdkyOl64whwkmQ8uXu3ptht89BtOdZBjIZe+Rot
KOCvVMFGtai8HhnrkKhr+HO+oLvbicfY6mNrYCU59VMUB5Nk6MaJWgxcEHXbnFUtadd+gnAmWY/k
NOaY0Uu5Ia4g0aIdg5PWboFiDZ3oTRk/kx9PiSijMmqSU8LRIbjii2iEoKqAkfic1WFHXDQVY5Wk
e8RWrpPNo9JFKtwDWDxV0Ep1yoSTqpudCu4JQrOKxIJMcENLYiyqncAdgpFsgVNADyqpUSNpLI1i
iOH6JglWUM53B5pDA7f5qFtTRlXVqRQa/BdnkSHD51nz9WaAEC/WgaMdpEHtxLrtIDA2lFtUcLH2
0t6ujq1PX6YpjxfIXSt75q0Lf+ITdtl4XfPKgY4i50f/+c4pBKoxw5a4l1bvRoeBfUrRRh3HtKJx
fXYIdgj+MEG9WtHYt3XFmdb4KguJRiH6osjzex0R19ndU5V8ShlzVp5Yj+Nsx+fWdhljNUjj8SnC
sZKsiX7C9Y32kD66+t2bHd9u1DmuHYu1XTpxToX3/SYlwLAGu9MBynPt0nuyWbkddYQ2a1O8S0Q+
FnEoHez/P3fI9x/HHZhpjtYJVeRMVfiwan2vRRVbq+Qmk97R/HisvFvgOvwVSaeXjJ50iCtITGWy
LM40RHJng6NkT6k+pGXpoMh7AAmFqI8Si1DPaaS6HfbZa1kcm11a2G/2MaacH9981RR7/yDr6mYs
ZjC95fBdMvewmQAyr6GHwj317N3mFjxKoPNCevqXU8qtXkir7VrOb1FgkAKhC+4OnjlJ1yPvG9yO
FSzi82D6utiMNKke/4givV8crhKhUTwxMaKm4SV7Qommp1cSkezFOYOhbS/o3wac8Dl1ZvgVd1NT
Hs3/UMuAl2slvEosCLPGgVTFRe4G10Mj4JMmYUYAADmxHw34QTaz6FdKe9hJYAzLc4ugKezfVEO6
m+hJlXvAWFawlNbpBTnPcThZ5FIIfGiJwl91fP2DVc0jd6Kn3Ix+AKDkHFyswZYSwFFKDtLbLgV8
PRAS/b/9wfgQVECT9dTyYU+VQ25DADRvb9L+C4GpMFFVCZFvZY8ysxI06vtH7j/dV2d2eZOcABXC
XiFpiof5sL1KYfvVzN51ghXnr+63NMXHEWl76K/2VxmLFBxQPGYYRTqGLRhxkzGISxgxJy283C5j
07nWP8qC34hTAGoJcx8x8x4crGvut1kK5U0ptBua4Lsn/quaisurk9gwsBK6IIEpB4iibgXU5pLA
X8KW6yB7nV/T+vlgBLeviXfRrkoqx9h6+7asglPbfiu+5YzO8h/GbzlqVjlimaHaE3wuCpd0Zx0e
6nLXL6Vkj8E0lzhBVqbXp7jJ5aLwYiLxtug+k5UOp+azOWRtBSJcn/maNrA4a4BVsQDVWU0cafqI
gJw1hm++D87oLteHsG3/SqysiwgmNkTAzb1VMaHuBUt/tnLKwfsLpoZDhGm7HtIdLX8h4/M4EgID
avPX1VVwHCsc82fVy2qM2rjXYL3+KAtLxYHuyjfW2nhE4uw8L0JDCA9Vre/72nucpl/8QWpf1fFV
4uQdic7wxooYMhf0J6xiJrEW5vEdVq/SycPnUMw4rTIKQNi9V6gPUNnU79bS5Wx++ojoqeHC1iOd
wwQi0zPqJPdmx0kvseEeKi/nJ35Y235IGcC54P6o+K8gYMCCnEZlqVqkMDJrLCIvc+eR3nhmbjHk
CKJ3DXCzRpB5/Ko6wfnoz5I4u6PjbyQHGxjiz2rvbo97qLaxn7lxhQjtphszZYh3LUQNDAteB2Bn
Vp9mz6N2eFL7US5yR8ckTe3/kmN6+QMLbl6AtrmSB3T6A+I9Bu3a0Pz+0oWPXmbYmJg7UqI1E4cV
lTjZlUF9WUyFHh9AhpjhmXix3oe5S8yJ4Ba+bkrHebi9nVhpqHoFc2IG3RRcUTxYAuFYInpuGtLH
vyVUJ79x7FV7Q072VkA9EQsAL0oZ6UgGd4w6JrSShwTWxEu69Dc2yQ9Sf/SGVC5OouYyho2Jlm28
DYlZs82ZoKS797wxTlrBHic7LYT3TuS/HVqolFo72zw+nNLdASeLYnsvZ2sn5Ln3NnHe5mH44B2t
vTQMS6zKi9p9zMhKoFuLYnpnu9FAzLsDmsqajg0tx4jZC7OB3rlWaYm7AwmyXdYXE4vgIhl1swuw
G94y1IZD7mW7Om3tnVpNGp6u193/yfgkzsTYeyfB92VyIKdpmG4zK5MIhVtJqidHs1DBppq3sD7v
p+x7m+6jqX6eAr35DmYrjnnGEHK774nDwr43/7ZAjiE39efhjrfYA5WnEl3abIPw19Kp7SFSrd3z
IRa7Kitd4iNJG9+4VwFJP2asRHPM2QmKwQHRtZMnx6N41DIx3a+5x6iDndt4l696v9WyLaMj5ppe
Z6ad/I8/3jo8CM21Q8skzKnx4GalApAe7/3rpEkyVlowHKJFw+TBpvYxPx22mS2fAy5gHe+r+TzM
t2MGiAHgVGOWldaMLoctNWhWUmHtqCHbD4M5IWG981CeLj0JnmpvOdZmK30JgshwLMi44C7qMSWb
DqUDtfMf1WUyWLVMWG6vrordEhdX7xVvtDhmKI9shapFwVDzyQRud0Jm6L+ZWj5V/ejFqlukbCK+
pCJjyARDe38zNepE3gloQAahzTqtnuIfc2mpbrx87nM3XilEa9X+etLcO0VVIzYjgGMFIplFYWon
mBqNt/JAtJB2QK9YkHM7Sqc6O4jEr2DQKMgoCp4+vmiw4gjzcLWdsO3FYU+Ca2zIroBaprmSby1G
2z0xaKtBoiN7/Ts1yPOxo5Gjs6n3DirGhqe3gSnas4tWXZUBPhhKtpnmGXAh+J+nyir2IOBwtxxW
E+DfRrRpVUQmMLAP5+DBhQ4s1efXd/D92WGjQz9h4F+ZXna40MilwJr/u/3rZOaPwVDl7kHayLeS
sz4hqHirTJSSQLK2YhxNYW55URDhRXUxU1xk84PDKq9aMGewIJjUXe0swCX5kedZ38WuAuk914PC
5Z7Dd9jeE1GhPwBx2oWSOpNw6i4dxgX8LDlQ6fzdPMjqvPWxvwyCV6xkZUBQ3eC7Bu3mnjmXyfRZ
Z0xYBqyTrXM9RbfQcZWA6sRKt5hxCJcqniWxeQSEYBSxlsUvsd3IHTo12tDu0SMOMgsCFKv01wed
IxytEyTtZICntxFKY0XeSNmkwz2BFXV+TAY+bJV9SH5o28VcIJk5pQU6SymOVXrk+/lobX2SRRQ+
qiP/s6dahlFZGwU/Kxz9/CC5APeLiRLLmC1xQRTPCKgSvA4R0RbC8P13uCifsciS1fu7tC387RUt
RoPHYF3CRNFviW2cbwvdv1854SEY7PqIl7OAu50jiFdLnmJrtYoWObJo5/MEv0N3Xjp5KhgNqzoy
LJeFHlajJA6Y2wcFxWFieFE5/drl7CD1Tf99CNRxVE+0mGrzolPD0DEILwYo23ReTibEUaFDmlk6
lpB0H1Tsz5OjulPAvhHUDvxDX40l9GSFrw4d+hgRlAMtotA9hNos+M70gEcA9VRC4tn9F983kEox
ek6E7+uTdLq9Luikmu5f9uXGYVJ2wjT2Hy8S+wsnmVa0F9cVjMPuKS707MylFsq66Xmo9F52JoxA
HwpuvWmea8r7KrMcQxHbOr7Zhf2faqAJ3XhNddxCYBMRGz3ZLAKr2rmJg+AYMXgIsCMYUHgoT3OC
JR4KBzjEn0n/dZN5T/tp4KcL/UEvEXlYnVoyzr6XA3n7YLzUzYoRPjomUhnNPR3DRHgT8vFfv+jH
6+gBdK2EemvmlHFVfH259L6ej1dtwDGvURCovX8hpg4dEndJy5J8hzblh3/YwfMl49jjRpJSpHpm
klTCeRMWrdQ0STUhDMUtlNYzNLErm8YQ5M7fAGTbx9xQDcgYAFgTFPoFAQhqcr1ECt1lCtqppLU8
Yon3K5M0kBBAsXtRpqA6RySSnu0FFnHdwB6eqG2iEG+uN66xiern2s6rlx3nyY0p9k9NLOaYLnKs
h2ITnP7/b7i333BbqfyQaQ7zXWdEv25dNBY4W/BVWb6puboCTIxRs7zg+99aMLuHzSp22QJMHMIi
HLgTa8PUnFcwbNIgI+NZI4Ip4wy1jiPVr8yh8U6zErJFWOBQiUYlZt3SYzkhWVDEejJynnlcclTk
Pvvc3cgNrWetEP8cUxsN4RihjjHv/Dr6kcE7VVb7U24Aa+se8CMB02ua0sXiRc2xRP61YtahmD8B
/kzq9sYCXMKHlCWzWCa2EhBB/LzpUQitZzOsdVMqed007wpFvvz50ZJEXzqxZ/naOCES5pzzTutv
6jJ/s5egEAGp/o/25UEUW9BDtY0dup9DvEV6g5YCZkMhTYQndSHTW2mEZWvH+3LjtqoOCsjd8aQK
lEw4nAcF3dtIEkmGXVnaco62MkI3IoX1Ew9h7jCkGYBIslMmG/NZTC3yvgHn/UDhOxESbAN9gn6X
IUE7AFG6J9aR9LmxxNnLVlxuj/tKukyFmG0PhSDOjEVBo6/HtVun+llw33ouzaNVXfCSYQSBkEZo
c867rhV/T6gIkedM65pbm+orHkvUx77VTpWdCmMS5E3N9SxyAiTeiHr7v0pXPCvVZ9I7HwtHxLO9
1zIlD/oZxGQKiLZKtmctrhKjS/xmXtABCL1HjdcuAm/hdEp0OD5FPcp2hXhCL4DxIUVgYulm2LPG
Yauc/+xgyHL/32djr7D6T0coSh2ZCUFJfRnCAgk3wkioVj+X7TR0bCxOS+1ZGNjk79qlhggN71fh
DXndiGcjibjSakm6ig80YPOotlDcp5/+xh5VMaRezMxiOXpK2gfFR4PELAJE+zr2oTGn4aaBNgt/
gCxfnTt1PlsPEPR89z/boL+gnbJUJwiHKsfv4ez+L895EqXqBRB+KsJ8CZKhS5sbcwysnrVL3+Rz
yaj0SlHG9HQWH4Wp2P4YxE70wzmDVlWfxxsEN4WNDmgcjPS/9U6vjdLJutFS3iDVwNTn7fx0d1RB
gnuPxRXeEIt4/fzOyIOD/0B5rOhZNBCsk5gfEHQ3OAylyEjHyohdu7yq4CYY78PvT2JY5ny1bRA1
Th8N+mJfYe32OURcHar/ekVWU0KUrLwqYmFfSKlMS+6qJWaOf01pejj/cSurfXP3Ho/Wl85t2jYR
ftlEuFDSbtEndQkpGecM6pj3tL0KPkvyI5OmNWR1ykDCJ0korA8hIonGbAvCComFCvZCUlnGeCpM
rtWeTnPkgiq1fA9/9Wq27eVQu8mmCwkXfINn+YRtfxeF4UcAZej2oyXQ2l1yCnjMJDa1p/pCO9tK
uL0WpR6ifMeOWsfwTaNsRPg6+yRII1EZjfci+PxXsuo/Ed3Tpr4mCUc0Y0AD3QhtbRe3m/h/qurk
JuPalThfYuKU9b54JJqN/91SXAieIhXVEF3OSbPHX7HBUKRLMJKsfTLFIiCKRLXlyi96XAOMP5dd
rt3QXBKQWt0VXRH01ReNdg/0gvSGb+sdTKqAxolZ5o6QmywhvrqGQ+zGHUer6BbbLaq+HzyANyHi
YN7X5bG7hz2K+22qu2akIu0SAfdTeoFfYZmgwcnwFsBeBDg/jK/r+gwH6s8RlBEJQNvL6NcQvy8l
Az7aAqaGeNqnIDlQRED596gC/8Sw+V/y09ocsiMWHOG8a3pmyLqOYOmPyYBlojqkAoACWCH8JeJU
9lbSXZTLnuWgzvt4Iuvjn6Yk7hyvQsDgEKpT3fiDspettBG58gSDVjDRMrtmji75L8XUqTHf3rmM
hBwNSXAKEnFGOTio+yyjJYDODntXcxsrxo8Ft7gilhbXOMsuQ0a3jiHDojMTopCj1Wun+EzWtKm/
uZFUWI0cumYRkxd79bLaiO7shP+BB9nFTmngB6qFH/AeFJiS41gAN+p3qC70thbjafdH05KNRcKl
+eMF/zquALm5eVW5WpzSDHn1JRcJv2icG4DxWDFexGiS1rDQrR50UaogQ4l/0PILkSKAU1SxauAf
qOKZeRUupJBwt0L+BiFU2fAaQNJlDAU3WZq/IJYtz4y/KJdW5jANJOGzI0ivpguf9JFLpRFMzvAp
QDXmhE9zc939B5gC22S+M2H6nDRm/7NSVqcvqk5zLa/BGVmuuXeLPnFcMPWliLrVMvBqi2CEfxgS
MAfWeLq5MFeo8HIdA66V6w+P/8ex7rOrTncFtDCmAKf69YoJlBGCtbwdYsis5SB0VZ5dLc7JNWV+
dwLpQnKqgh2tuCj8eQWIxYELhRB+OXm1bGZJM4VNk8c5WdtO/hAwxbwUBdykxGXTz7YYGhqXG5W2
2NJJ+Y1CDBFPHAgksbUCXCo2OmGIuPdKuwSr1mb28htbAqqJkZs6xdgVoXJxflcu6LiIIzFf3RN6
IJSF1L11fb7GBZWDG8ApWmYXLtgONNdivo1OvD7O2bLEZ59blET2uNAJut0TJp+2w9Pr4JjpJ1h4
HBWWExBDRNd7DGOFjTum6wgCyarOcJ6gcknbwAcDRbfy5gMMTgI1kjNykffzJHl/F3/pyYoJtzZE
bShh8Zz82vSS5yKVh7OBzXLCxu3Mg8HfMDvhDv9wX3LOlVobxyH9XmnX0rp8FtTWAXGP2oeMFSI/
TXAH0qGG6c8j/FNB7Do/9ry2Ae5vmMd7jsixwcT+AO/3psg6X57+mppWRrG1KatnZrFcAWRuP/wC
G+YsnRxtdXYYZ0Y4yCPEE5DfojXcTTrHGUSAgMrRlKbFctYwJIGQalGC1QpmdF6Pf1x1p9tE1ZMZ
jOkn31Q9SyBTTua7FR+Cvm04xtWk3vCuKQFSB1g+WHzs9eK8Oncr3pxw4w+BjYtZXJKduqhUmWqj
5rxfehmb8fDD5IXOVVeSEjLCtoT4K5tCUseXeRPY6GY579t650pwlK5lIScKyTNg8yiMU13Od+B2
Pkq4pfBZ21ujOhBIqd3oG5db1Yj9Ab6mF+E1LLmH7q/9obaoWoICfdp3UvAzETPIpELWGAFjJra5
YscfGBU4K3BdObJHq/hJtlvPLJJWhxpOmQI8waRBGDQPfE8rN1KZNjd71u4BKp9mOrftC/AVGliL
FHwwJuXEfHkkowXjz81CRhVC0lYrxtSsFwCPuH4mnTY7JSyoz1c0882m/ESCLh0RiCJawZuP5vXj
ykLD6W4dS2KIkuY9SOSWocWXdmD+HIEr+MkchEiigOxiGNvtsSZNmf9jqNjbCPDGm8u8pJNE1ONy
+gKBZ7lSeg7mZq+Tw6z7NGK7V4wY2zKsOjTz8s+hDTMtUM7xhYKxwsechI7eV2SdZdjCl91esyC8
m+HT5RKk5QewVtldvF1hAz+lOQNa/bAwl9sXo2ASuFXnwQEE81wReuIF1XJWwClbgC+5nG5LlQ4Q
ob9Q9YHqWrHVXvjPA9YBFvSKmF/3TUYJY0Sfn0Wub/PtXd6A2Vxlojj1LWG4SaayyN0Fz3rc3zOa
k809+0No7WuFE3JReMc3uebrh61OQUWdRyL/UvNPpPij9gFTpVms5sVYsnEhV6YAfkRET3NOH8CK
r6fd3gvXLYSzI/wef1QhpNccbDsCv8eTPzePKIyYbHipHdNtwOp7GEBpsMPQlkh+VpJO+uMaxoSI
qwXUkLn+y79uOJklMOjCLhckUoxF+7qAKyDqSGpR99AZ1IPBDLkZjN2XrU/6zD2dUnktaa5QHu68
Zfr50RMBkF2njk/oBkQr3unc8kzNK58DmExdTk7dXEVaYD+xare5YcRUJsO3aV+/Xqpzm6K/bIjv
AG+7HoXgs9pm9IXB2Tl8eEPmlIonUnkgGYVvuMOo0SgqudDU9GRtvA5jGjsWI8hkBrsHTsXB9Gwd
lSLUu7SKlyv224SgDoquv9pB3rryxmYbzk9sujeD0AfdNIjRsenRnA+qkedr85ZQ4WCeFi/xVWst
CndW99cU851/4t1A/EacPddBCWv03A+rchSiEFznYWTF+Gtl/PIdT0vKymwWkC/DCb4Lk8O7cYlC
JrKfC3C91Wn5KhkW0zlLQVNcHwt64Fxw7RqbgaVm8dlk6ub1WiaaBuDuMs14go7uvUz2gRx06Rs4
83uviDSCHHLLNRq26qb+pkF1plLBv2+KJHrK7fipqgLxDA5E5S/rxUy/NTpr9rrDuFfLM49Sx6so
DS15lyTVA4Yu8Jk8imnkbPCnkihXUet3lW43okOiEuG1GxVWaTIANBIOhuFTmkY0IGwnkAjmxPLI
M0eyYBWyVTiLetzomcUwWiYGOA7IPBkGZFVNDTrIjUm38IOIWgwX7YXORUWzwjFM2SNcSDGakIBM
uR6ywhHV6JePSlxL3QKPYGuDXHu3+1puQnWKM8WDW5p4zHnEPJO3jWWsFk+5XQbhE3X/ODag3eYL
lEGUNV7rkjT6c0ZhGTLOVTRBmWqdi0WO+vQ0BUFBVwaI8ZaTn3zoigDGYgjUfUQQrV1WBiiAp4ee
EpZ/v1Wb7ngeTD3yrK3eUGS+CiIQ3F9+MhH+sYSunv42o79OPbf61yd0bjpdkJBy9KuNmIgZlmoC
/VwDYAXLBeTDKAr9UqurKrtkGrFtVJ/Jcv6GS+hEquAA1DDLVxncvY3ZwntuMvCtYTSnTvZ0yEwH
uCVUWwhreO323djHX3ffInWiS4sAm/YUKwVEhg+Nd5ud9ZBSEf39HzHIHWzqolE/gB/rTjhh/oMZ
mfWCrIdf8hDRWnnvgfjs0dU1oX+5BS6nAWuZB8ntMQIq7ksIDNH/7HoChMSCAvV6LARcMLko611a
CkipnG27HHXLpGX6Fe2Zd8VmT8hmwIAOuL/Pxi7jKD7Kyi4dmVhOcgNDxkWggdh5Jh8a2gU2qqmC
CwbBVTSGxR5RFX2TcY7S7tdBzL8t7Gat9i6FGarH2c9o0zJh0c0TqzKPgKljnCx6L89zYMGVlpbu
QRSJQHj3lRvk/8UB/NDXBbrH48VHPBs+PsxjFUIdCbljJI0ox6Rx2HrOOp04e+aGrMNFWLI26UYx
tz+C2r1PFdAnX3CQsc6kCxsdh0ZKF353ME71AcKKlphsNvSRh5vxiUoJDYzPW6X128hezslz1Edu
9TiNzqFNKWBGAGWr4JQLH0qydG4JpxRJrjJRZXnXHFRA/ECYfdPISFzF91nFMFn7uCMp3p4x/q29
oM32pQOjcegjpsFEUoBb1G/DiNNRqAAA5oPTDnkSRxsSM3AWbQAkWSPaS2AF4DYLjiuVpuyeWgEr
puwdIDAC11WZFPsgtXbzUrNwlJsPBnPAYWF+tpNvqMb5Ch6OXT4nSyLH/lYZUgF+LolS4AwdC4pU
m5TacYSf4cHU9UhYqxftie3ANlWTu/1P/a+tNlh7blT5ihB6X4UTAxYbJofE46nDvOYDSq323jqb
x1ChRIy4laaojVCXxy2f5xEFVsXWv212n4HvIoii05BgNwu9h/4j2tPy4UIdYD4e7GVtahbWkLML
JqY3SsUYcaCBGaOkeUVux4NV6NxP1yNDabR2zivzbxOhultb4HdveRbAtaD75AieUGq3xktV0J5X
s/1r3b4T5r7JwRATSRHVZv47mWkoNBfK2oWV/aCOqS7rAZcv9d6b6MB1s003/MjUpik9Wat8rPHy
XyejbDhVetTRvtrWzhoHVrPjydXZb9rDoH28EmkN9QHH/XmbAS6z7kKilscOzcJGexnBULHCNLJL
c/kByK69E5RBbuq8SqsGH9XfwS+wCtqfwt1UH6bz6V44L2zdNpjEfLekNQ+HYR95lw5aeHo2BlFk
AOqY81PD+TqlI3MC2ci3qefC4ZvVEYu3/uQYoD2LiAVyWwrfJwx/7vEPmHvHSWWzbB+qg6p/8rVs
qhqQebnf8FnYA1U1j3nXvZYgA0C4kJtrHPyVKs772ZdgdT5QcSM0lEZfeIjjy9mUUhqPaGCdxGZ5
0p1r7L5rMYN3Q3LX+1uLHpvtKQzQPiqNfE6K31bfXD8jT517AdzL6420FZ8/9YOy0L5AMPPfeFKM
hqc2FJp0BMqHkl24s+H+X8yAvivCiK3fjutpI7xIK9L+0nql0KJeQ8+L5Fpvv9TaOV7dfW+YD7wO
1B9lbRotKlWQkeiZF5GdPHHMK6dxLH1RP/zPPRr5DS7wsaM16s5/nm4tLTn5LINXD+gCU9cjj+w4
Y7x76chloK81pZDo4XhxHZhKCY0WzU/N8ozvEWLuhMWvS5H2rlyuAIAT3w5HmRBl3VOm+yODabrf
PqBTJcyGqBfgFba5a3BuRz8TB7ff2fBg9+zXn9bZ9Ma+sAhQ02m0Ly6labH1bTYARdO9357aMrAP
Hjna7/cDwsUbIKK6R3xhRKEdzfUSvzjKMoDlQf1DZwogzDrwuBkU7d/yWpz1hp4u+aeNetQ6RWTU
N/fZ2kw5X4/YkmEJaN1Pnnn32t+P286WFR9+1gUiwIyUMXgHJpz2aknlOkq5FkCvdpVy9cpVxtd+
BqOS6m7GRXr6Qw/ooN/V9p6xmBSln9jo2sKqhZbtMFiKghfPh6MsCbMxKGAmf6one/uZarS6SVNW
p8JN41SINvgAJGKKIKfBq4FO0GiBLiKw0IJYbQwDr8HXfThCfWPhZJt+xWDgPxxkhcsmhOlXmhua
zsvbucC+LoYZPbKAk929LhPp/Kym+Jfxgt3xTZwrESmhxTVpesOvWvATmp7nZKDmIY2WySSluSB1
BAdGgczpGJydSp8ugRbLf298kIQNBBXRUA6Kqgy+WdhyScXca16V3s44rmsboK5lMUj4I36h3+Zk
AJJrwNQy3yHafLTf+xOSG2n2K4D9FUeJkQvF1JQkKXH2M8YodWz7jGA4WMbvsKeN3AnMFantX6pi
lddKMXv7wJgJk2i0K4jyCDy0hI+X0n+fPPDvyU6XwFb5v3VcDND2usopmH/yFuxGJ+JhT+Dbm1Og
BtHQXmO9GVqzdBffhHZ4X868x6ENHoEFN4kHaWyD49jFfAREit6GHkubq8V9ZTL3dDZFUZqhtRJ2
LNgh2zVP5mpmO6x5/3fAM32xFBuRLzKT13WeXmTKbU3uLVhbNbXCoCesd1dOdbjZ4Zp6ypBqnN7h
ex8+8SCikjIPE+ILWAgtCGtwn0i9+dezq3szVV05S0bZH4cwG8reo+8mVyqIs4V8DB3qmbHjnD4o
GM6ExtJLPW5QoL+uOgDmRrcKWZahunlL3pFQdfwv/pgwCWAkr4iyYm22GOLMx/4nZW2yAfTkmY/N
w80XRE0EWbZM2uJ0NY2feXeeinlH44pIH9OvFblAA4i71dMAREx8SNNetU7h+IYbW677ooxWkT8I
gqGTS2AtQQVRVeQp61SaRDFYLct6BimYVIAXW4skBs2vo/iDWiu0X8p4XvvLdvmLk2opQ+Zw8JQ5
NuuGfUvDqnmZSXpsGp95pSfteBHoSkQyi7688M1PUMN4VH/8QCRY+Yf0jgFo7luGT0WgCzvknmWt
Pyp3cMwK7yx3MX/7s6Jg11cgchhnjUjg0IDM4vMsClBoW5eZdKilu6ZGixBo8FDVGYPFBoREqGmk
31LBazCpZXxtAnrIMD399xAORArEZFgGExo/JTyrHlKeKwGlFKiMowjJO/cPYiIRnNfANXwQVMez
NBebA8ftFrMkgfF8/sZfpnuzA766HFjTJXarsFtcHfU2yxkhg5mXJ4Ydg0ITC/GsNbLxeAHLz7mS
b5bRokizUPhipwCDMZ3PclooXepEqeBvNK12RcT3azUPOeOC5d4IYQLwGG2J8/WB1hYsMGi3q4wR
ZQ7UeRaHI2IXmXu0zKma1ZRt4AxrCtNwfE7aRYHpZhRtgq7Bm8aXlmjGHCCEquSBHg5oTmKJuRa9
5O9Ujvw6O9urYTvIJzeUfdWsBXvruWh6+2FZPLfrAgh/DNUFTTKRBwVbQ2/HR8kSm16F5v+z2xwa
jemVzL9302LG2v5eNMLO6DRUaQVlonOMPeuE5n+gzdihMkAJYx79ShnWfAaFzmQ+by1kvf6JJpVo
XxP8U8oHXZfkEQlKO0vjP0cfS2SbBEqXowZuIkg8GwQXVIM9I0ekwEG7ZqCE1sUKf2kY0bhbWMbB
E83s/wAP9lRTpNW5OOn+eVWfCvy+byix5QQaozVHMHgGmgCTLFAELivKxq2cDAaZR8tpagLt7s57
vwzTjxPSr/3r719KRycKaaPHC++/QCL5Et8k+6RW3AhyhQviAmGPKA2FguKj+97hwX10KfndzOM8
Q462QmVpwuG15UFxHysx915Xd+At+7g63K/cblby+8CMlawYSdSENHzXSM2+ATA3tB8qapMgcv1k
JdrA/N8CTzwKyNItoWR2CuQ/AqB8jOEipD0W9APLakB+CbnsRDe2hMQ3ZLCIukuPe/QG7qF3klQH
PMYpt7pxAtu7z3vB3EPpWe+WhrblDh/YyNxg1FPawrGVvEbf6DxU/AGDKhSAC3dpOWgaoyFXb1sL
9hEn+2yNSQMnZnw2QwH4xxd5SoiLQ9zbAfFbzW1e3LsQGVuAwSS2HPg/ZpvB/KQ53/b06aDQuBTs
aYSAnBcAdTILRVLwV1PDPhbz41l1pG0/nXZ2AveI6v5qeL59drWfwY2OxN0wnX0MvvahBR//p2UQ
B3kjV0Vzion7q7d4LW4aqMzoxFShZmtBmXdAOqEz+GtrO7iVfzNmcpvDiAMmWZ5Dm2aS3joguAzc
8/vHuubFcOOww0aF4aTcNiaxrFHSCe9fddlWjITJPWm3vPAEnVDb/VXqVSaN7u7BaW74ymdVPCs+
Rf2D49aWxYR0GFiAjv2Qrbue7ehy+3Jiz7FIf9EMsBe6Od4NsgetKYmsZRE2TFLNqgtYxJWw31n8
aU7FW0tylMUosbl9GuVO9PYWt16rMPd8QlYXclZ1VY9uUfgOJJmCewEqrA/KVCkQcf96sZ383ZGY
ku3fbjM6xB2XFJBALiYR1IIh666dg8oEj/HOBi0kMrJLOPbZr44UDmDG3mBLl1YFH3YruqzBDALL
8GsVbZQjE1Ch4hNsihuWiZMmOhRFvC6cpIdGc83lXKabApKjAHz8hNenaztbxH3X/Fz++baOjW3T
8RndbZZ8ekAod58jLU+zLP/BzlyqKfAxCPhqqY2hmXs1AQaL5eqXodGwFeavm65YPoQe/btB2pjC
ZFzNr4/hvbOa73Dmlk3ScijZI9Ob7K4qqmHeHOEuWHSMJoB0FKnckauSJz9Q3qWkZA/0aiE22bmy
1SyLyzwQ3IuomsO48TV+m9uMRCq08yOotoh3za8bUawgxpaWafqZNYjv45/nn+cMFfoTWl+4GPjG
F9j/MIgG62KVnxKAO+4InJhJgh74kThPN0E64b7AC8n9FZ7HH8Ls+h5cA7ciZ48cj4KhQuy84O5Y
lyWXFAOTpKrXq4Gedasv94hmNtdOM/r7Vdsyk5+TNq2l92IIUPzvvha4I+T9vmG6k7vaVFmMDRxK
2b1VYE7I4QpRJsvyCZJ8B9v79glh4hL44F+JQbXsJfpfYWg8Wndw/IEmASUKA82ktVd0jwBuh6Wn
VmJUwvv2pqGENVfvcHNfqpMCMh0sN2S+oh6ntBWaw7KIWVHglWWvgmNm2zOd86UDn+W+4NeIBZa5
/fIpgeM9TlGeTqns7QyvnONbgATNZEZKhjqbp+orHjlFO6qQ6shvaYlbASwJqS6Gvi3dDgN17MAY
GhRRfW4SOK9sWi/Ofu+Fiy03Rr0UsO+R7xtVGvmSq07WXrSfl0AM43P6p9UqfED5Ec+ZQm2S0OeV
zUXPZ10tCGsM//LU9RcCbtukhmssmL1Drf8w5IymfLEKPOoQ2xL3dckmNy1UPJVzP8WWBeggMJFk
tK1eBobC247gEozmdLNV4ghjAgb6Y51p1F/2hdQeSifhR6F0fQdMO8eXrSXrs5Ao3I7geRJeHH8a
1mIyYi7quQC+ClyNvTKyLj4XoT1CorEr7ui8DoDkt38IvO1RjEI0UsU6OiE1xtcxsAYb5vG+cx7R
CTq/tvpN3LKDUsKZfJrPTIIj9tzizFg+8xZONKeMrMLipSdhIqARzzBrPbmIwU4SDAYhcfTYcg4T
9kWFb3tj0cJ7bjaiUlNnF5SdtLadAYRic+831X+L/kgi4kEGc9QRTBJC+yJfD6yIi5KmMOpJiTQB
Q51VMIHJDkPWSIgJMCP+/CGI5KVMPDgNH4BPYNzrtLhMdM9gc0Tz5RckFuqmAz2ubrCYg1z68JUv
siZYsUnKU8m0qCOtMoTBWdl0IsMKsZdrJ19nH6B49iBFn6LP2rvVRTERjoBfXz0BL7xnId1SpcEd
nJb+MgLnJd7CWsWOoUt4bwbhEo6lX6QEc+eOPK/mfcuNps/BG3hNNevt/C/tgof0F1nG89GydvF5
wuanoKG8qgoU440Qqox0syYayVeH+dMXddTZbwxHnft9+If/e8J26zZUS9gAjc6gDXHBIDwJ0Cxg
sYzFCS1ena4A9vbVVJybDuB6hUYZxDbQcOotOi+KIJw/qffYRODuAGILC+lBHAuAFSwicMoHBisW
DM0B7WQYRc4mlGkxNUAfJ8rtFzA84ln3rKCAOMXqAe1tzSxMhXn0sVNrHY6WElxnliNgr9x4K9w4
TdMou956Fj2GtegE0Zh5mikxu7h6meDaQOTaQEC6f9Y0R4NKPhScuF4thiJm0ZYRWNBxdJUw/Cew
uJ3eTQCkKsh7UrMrzCWiU34gqMKP9uijKQo7HpM+MQP4HKuVkpmWBUVW++o+KmEiXGAnh6LknNDL
/LkXZw4qhdZuw3CEHuKgxdPlL+JSnk8cd+mKcnxxkd2yPNOMNVwqOJhO14hGTZrl+o1lZ5WPNOrB
fAcmbCy4M5EBho1JCBT2fLaNU+GRLMus7EucjS18fp3GbKMou72P2vv4mrLIUNh8e4+jBUuAAH4s
37H+/4M7qfZgOTTZdin+JMqAWYO3xJFMyBubUpUjkusZ/ZZakLEXnkELkuoySR16Hy6bCtKblaWc
pxUjjLFqC2dQdU6424z+ONCCZ+8YhtN+ew458b7BCYqlhgAFlIXuRqsYtCAPhDcLt+VuYN6l7ami
HS/ICqbGY9tKbed3XyRhPxE1EwwMhG20xdK0zgyZltOxDaX/SNqtCV+Acy+kFlNQOp1sFumk40L5
3NtzGDAmkuTb5SzpfIjb0m+bypTDqATEY3YzDXhbEjd/gObtC9qprSr+bRDrBNUza4yOFzJcnkFX
DmYCWJfkwEgA82zEixvVXk7GtwvhxFVfc8XkVXySaK6kaUZurfdzUcWh1gNJH7Lr0YQET0g8acRm
X7b674lBQ9IDUfzTt6ujbkt1e/C0PUWikdYdME27GlM4oB+TB/rdBVFt4Aw8VPezU4Ak0xxI0t4S
F+ZH3dAB8wAX9a6NyckwpYjjwbUc6gwn60SU4W3uIrjobfC0H3ZXp/DqPybek8pIGkpABpEJFPOt
1U0obZyL2Ulo3LZ2nrbQPpZIi1n/ucYdslrSpWRvCDS33nAW4GdvP5eX8m23dAjSW1O/Vw3gGZ1j
SSMh9neRFZIi0sacG3kndUaWeQbT+ztFFl9EAjYvl8BcABnmSowhUnEAMs54IuWk4N0TqH2iCXc8
lv6vPWyq7qaunIf1d7UE+3OFDTIE0DaZXIMIOC75IR4pWoiw7u0ixKQ9TekvYby7VoSbflhK4qkY
LRJ/Ea70TPsEs8oU6ohlMjqqFFQtXex9Jy7Gb4dSRpScrkvuTqJLjxCpjKosA9j7DLlSlw9XpD7a
SSQsvYmkjFWK5OUE1hDTIjgHU8dcW708rVKKBhhVNinJGJG6kG1tgcqUZIdboOCl+tAVd1273l3V
CTiLDhzy7TkBVcjNBAI4dthRZTlWcDpqqzM3L5E3hpk79JRltylATLWlf8Ncfauik7l9SIzyZAnj
LcBSNEo8fuoprXO/QWqdcMYThsQBf42S9NfHFg8hTz9p0f5iV29NYeh9/gLXTYcuOw27LhyRkUoI
vUAy7hxHlTaLH/k0U3c5j9kahC7muKSX5y5wkkaIgCvnRtXo+0oOghNhuDJCnRO8h/UzS0XGCOYb
cCYnWjkgF4BH1hS/AuA4M+0NQt34ZSM+fEMIcaRwmQEESMxhLQ/lRcyCqnhyq1U7FCcqjQH9Q7TM
MUJIQxJUDkqViNGSp8Aupk5sG82iPelreJMiQ271FzLJ5S949Sc4lHAzvdavyMT/XgmD8Cn7QsuT
7SnCKUetvf7LOhn4CyGB/n8x54+btBsyC+7+/3maOHzjUvDV1lfhIoLF76Uyd6HVWCUTLgyEbRtA
dye9eJqJS+FtfWu/TQmoqKx1tTzS1GNhmojJG147yBsT8nushyDrSxcUL2O7cDNgkeLtcOPYKfRD
ZarzgPNKupbvLc71h4gzUQH7n2DTOUjkvIdJE1Aaz6HpoGCOzYRgNUXcYPes0hmdhcyylF3uYiw7
YeHCfclO9DkoGmo3/lG9By1xq+pCzf3SXDTUmSF+RK6oX9opZ27k78dltPXO8ja9LufQ68TGLhTH
f6xX4/wt62rGDYyl5ZQ5JI3ZglxRjPlVWZYd3CxvDhLIrYEzUmNmS1mOgTmj0cwWxsdPKiSZ2hna
PkuDUQzA2fznS1MdPcikr1jK/NKnxD9hnF2erieTfT2z3wSmyNWu3tDmtqFZM3sjenlFNDDLezAO
TrP+HJK91tojlTlpZtSDdomUbALDB0FK7uNnpHw/DbXt+GAk1jLTmw369wk6BFBeJ46msdTtdp+S
8w4L3Vv8ryETv39d+Ls54NAk8YRtWAAEIM7UB50BdIu3nbaG6OUlNgZzey1fFeAYpeLWyFJtNBDS
EcY1Tpqq3Q8P5OT/eWHjEfnFPoztWqqrvR/z1tt8mYwLRwXVznTmrN60qQ2kh0Y9r+UZqg7BVHgQ
KUQg7n9zHQohAId7LtZGYfyc9qigAEbhPmxM9T1Y+CiUyaaluxlyTyg+VArYkacrcC2y2D7KVt/S
rtlG6E0aL32APXpYm8OMAgvl+mpexNPq+q7t8cet15EZsnd2DIh1gr3AGJOmcfy0uni5exUG2BAl
+yRfpblQt/TEwm2lJKnr9Q75uDwynktJKbdKwATuvU7YB8l3HZa6rqLzDg8y/g5BWaFYEd5go3ko
xo6mM7KeMLdItDtCWm9gW55dpZZrPeTR5dtuzYDlLI5siZjBd52D7BkDM/jWl8kMg21UjkYL4S3U
EjxvmAXwy9vn+VSL/4yEDJxXfnvjKWmtGsBEKkWE6JVVHEuDIXuBZ9T0Cdlmxlqoj1BKcydo1aoS
pKSPCtnRqOJ6xO80QVaP/i/6v2DRGBeFeanM7eCwnYi4fi+tW18XBvbk1IDsptpZ6Y33jl4EadTI
bDQ3qxcgt2ZqV+ggQOa2apuSqoro5u59sOKYWH5Lsf70HO73ApXkeq/hM07jMM6t1idjeugUJqP0
lfDiyRnoLEvJrqPt2V/RVbSPlNB/oNodAn9EGbBN7sxODQf60kr5JUfuISztkkhoaAgrzMVCtWkf
W6hE2ZLBzbFtG6FxGEdjXHzCKGBHBOXk5viuERSeFvTsvB3PHRZLiNcCDby8Sm2Si7ToL/YeaLUb
cQgEF+7UE+HwIwRElcPQNQeVhAPlGnwiwEUIqUKp9WR7wJ3DYpqn5+KxxIvjNDej8QnqlN7o/+u3
l89jGCG4bzWttJeZ9RGphEsPsuBE9Fym4RvDccNCdR0zeGDKNOyjDUdsiCpgPw2zvbI2uAKpuPQ9
vi2DdKnGWxx/uJPp+OkAloA0lKJnN2xsn/v8+n2fm1Zp6IqysMkDAeFTJotWO4ABln9qBJ7Wsij/
I+FJsCaMyAQvUxYia7+4M9HNLyfgIKrDDEeFCU/pVNiReL0zrqP+GB5lEx47mleiHNd2PGD0avZo
OTEVTQq0iTJgnPyQ4KKOa7JeMLQpi8S0BHp88vtg+9mOZEhJ3BBjneyhFsy/u37rkMh/WXP6evgI
67TaBPgUMQnmkPILd5H2gWXD/4XWsGCG0EmfkSdPGgYqZdWBIv9okNpOPO1ZN0ZvxBn5km991VRk
dPWxXeE04TfkZWO4pA1oKvjoVyqmYB1BNcQqbL7/BTxYioEVbmPESIFRWWf3a53rYnrbn6sAftFd
puzpd3RVB1W1feex7xy3OtrDSkrocO8ZeaDcQQQf/ycR7ZM8kfXZ/FbXUIz33MVUfmCFYDuCTux4
b6J+JhaluLWU8dwyNv0dL2OVpYJ6bBNlMGb3c7fB69+r2H7rZpLXZX5g/T9SP9LhIPGwYSeRt5Kf
7G8fzaPVxgjrz+bK++ekhFSFzPXGByc7oJ4eunFuePPs978HPuMrTCiE5h3H+Tw7Z4fKiHMvkVnK
P4OmayubosYgPPM6cK+OXZfL3jFmD18BxAaJil4GNoSMgy8c3gDdNdIsjrwcTf3cjrEuLp+GGPC5
l8QFOJ6ktCP0ZoYFbRjO4l4Xk+9w2QB+oiTS7voZ5avlnU58Xm215EXzuCX5RoIMsArvkTsAETH1
BZ9RO1CY7Sb4j9/zWLrrv7eAMaoQP2OtYlBF+KCxxlqQVk47SReNA1rrZaCi5ohG3y2v6K2ajjOO
l/jtIr24p50FzY/dZSLZorNDgoxaH/9b65S2ariSKgCzI8R9Z7gKjZTkksQOOdyFHm1SVJEla7t2
kzx2I+l2vPpc7nRLsiFHbMLdIac8rX98J2Qsw/ROo5U5kor6S/OwydFiFBbG3p8iJgbClvJOOEuS
acmcnTHArbPVPbgFMrCWwnF/IoKwPH2yllIEW+B055IbkAXpGwYBbq9UMoMTZxJnWCdWdBy/QtBU
SYW/jvYEHLSNd1RUdxP+kzTNpzWeOU9uGSYBo7NH5cqDnUnwLZo0EYsIPb34QAICQ6hGhJJsprHe
tn7A9Z8tx+pojacAkOJ7lFouhvGA7RYzRmIpJPbRvouxu1SfP87aJDr947y3A5vSkff+we6GoHuw
Wbw/FOp8yrXJJKqGRMdd1QVI/6Df+rRrg99CBZeJXD2u1mOp2dL9JAqT2/9cI3blUMJ9+vGjNd9b
l/7INrKhooimrGwragscyLaFkZ+Y/jyku73ep7JPA8q3YFuPQaohQvTKQy+DpzNUzrmIPJJE3XjD
ik5MEaW+WEUCxNOx8FdBLJ4JQPDpTgg/k4KIHGh2Q6ofDCm0hNS7x7mJ6YEB5IvYDLtG3UgSf3oN
ujzJ2xPSY40MEHd151ppXlUdQ+BLzk2AQuc8L0rCRzxHIUf/9OETrRj4BR8Eks3fHZhosM7YdfZf
+QqJ2rWeYw5QGZ1ffIfLiGojpEQufJF216MjAOP3LY2Y1fTDjMrATGmY5RqWEOZyVjVgTViuYVhO
PC25eQ4W2mF5jbXiZeZ4+Ee6GBpZGjT+I53ppPEJaz13WSAYPKBa54lzp4OdNsC+WagUL9KWFjU6
KXTZQrfHdXBWlgCXectdbQInMp9wtd9OOOxO/upKnv+97MMPFj6xv9CcOx9Yt7Qpd17REtonL6bC
eJO2j2SuwOmFHpaOebToSNKzKOPkxjZvnhGmP1O3EPr5IJ62d90xk6D/EsOqfQC8SUQ+JxI8SRw0
MPzBVgWQC8Zz1H378Q2G9UM3hKSVp4nlyqzcHokho3zm0YTDf6eepfldWy3UDRXMp0dnerHdFkux
xaeYzq+uR6cLvPrB+Es5LS+NodRK4tiZ+JenGfwzKyiyUN+KoGwulEXsDSUERhLRWfYYGLoIGKLo
KnB+9MDIvz5L0fwFx9wdUDlSrx2pMzHIU0yYor+wDQOMcBFkUnZc4o5gpic7ijKvT00nQEPw63XV
SpvWBHFEHeDxDlStuiVPzi/8CYi26vssaCMfny8Dw/zjDe9M2xcogx9wy2STpRsjaNZIbKetvZVp
VaP/tE88ECePplg0sm5gdh4cYXJ7l0Dj8/Bm4H11yu6u4JJyOctAWUYRn2tOXRqG/xCXC5AePEzP
a5A6zT5aydD1+Y7xJJ0YOaJyupiubhIso3AdJAxwDRjsW7LQ2S2e1u1wM2k838Psh/AabgHm6Mal
HLIY7rlBqye26e5SbPbrASM/ZQdl794ZZqb7IBAyZ4xe6yVTMjd24Bg3Fl2slrlk6oQ9bA3oAo8E
O7f0umyJLjsIFLsK9NgvgSV6LgodqZQjbZ+hKquCNgChYDAopNrE1icXrZ0lmsx0pqD/1uo87yvo
Ac06fhDcxNc+J9XdpKrzcaPu3zy/Kla4q26997LVqlXv1cmAfpvZTIyAk8YyjgMEnWxY3CbAMpvJ
41uyQByZmLyM0dUzlFnnl2+j8SSLHEkkKAMqXAOLH/XubW1oYeZKo0QucjTO9rPHveMCSINZ1umG
cw1Ax8/KqCTSS2ByX27I5CgKCkC87i1k2M0HcxoqA78SruMDgEHbqf9tSc5qFHLcfTdVmVUzvcjG
0pPhEQeAxw0A978lKGo30eobER+XycEgtxn/RsxKaXt+TXalDXod3i6u4HVxTlhQDcvjz66UrKUa
CYp9cuethAaIrGgoHTQuOoPd74VsgdSrAH5RkPiMTlKgIcw5SkLbdr8RXVsTwy0oWkkvaVqwkzBA
TUl4wTdXukXSEGiCDUaJqUoArS+BIU1DNmOYJnB72DLykN3v9ktOz25bsYPf0+5Ogh9+8dGgTymR
PbRBOBdxQ4TXWV9iqNmxsOibvf2/1awXFjADeoFwfbmBmlNrlgyUOvPQHmwCm3kBmRwoJrauzYfU
X6sp4jaEch3i3b/UDdqdB5MT7TNRNPQwmmCo7nO3FDGSvrmNRzcTFtMns354pO9EbhmileZqrsRp
rBiQs1K3fpxxQ/mhiUVBlR7BkBwS9EfuYMhKXzbS0IrQJXabu3NYkEHNOEE37Mx8lKkinDa6DiSm
h74VLP/bM8N2p1zE1SMN9IbcbQKPT3/yuPdoPNSJfoiBfrhFbhnP+1Lmv3ycAWelR5vnqAFLTLLo
Br2NDaU9GfMF0K39y1GmOJFWPLXQb75SMOQIDuV/HVLbNf6pOATiI/oZKLOSxnQPF12IN/C4qb5U
cjGNjFDDo2zhYHv/42uLEMTlFeuX97ivetkSB3WUyoS9y91mV3sGnsvV577flpBaN0KO7otOAxeY
WOG4r5gtM7PZMO0E+yCDvzlp762GQsESF2FKnbL9L1jTys6NH+8eBeTyCBsYDKLtnWDE0qJRTzbQ
ZmLa9Za9FisJJ61X7HpjSL7vyty6eU1Vp5ClZxUDHDIFFaIK2sjl9gYkAEEU7xkZg8PZ1VW0Scrn
1fVpapxAJNWknpAxeDLa5IAJktUDZaUq62PJKzgHxd1BjtNtZdJ+L+JUPZF+QhOx6Ay3NcpjzJ41
mYlHUErxasSHbNQVBVjcSRW6tvZBfG5GqpGLO0tq9Gk8gq2Zf7rpfLEUC0bOsxFyMcFgdLNK/Z+8
jC7gNwF9EggCDoxkfTXIlelcwOUMBBtSacqVP5WtIeiLH9pG+61s7k6N9dPmm23yi6qLvvg83pBE
ByzR9//oBpxPDpQmDqpkvyfXJS227dCHzGM/5XDVlYf1kqanYCVNdLUHwy9KB3SgDdZ3Mz0J1tGU
scVPZStBF01c1m9uiIhcPBrNDWgBVLtANrBGKSSGLEOnolEBgMdvbn3NDwVftYphipkV8o0GsUD7
hiPLS8ExGt4fA7aEW6L0vR8RZvxUPzT/Z19D25PcgmETF+ZtoIX+5Qu+zrkxVrRmeAatMDK2pncA
M93rkf5lnLJ9Wyt3+cLkR8ya2p2v4xB9rJBxpR+nNTSIVoxzMNJGd1aNxIDKtTKicikP61vbTM1j
VKO224Vz+2R/ElkUOC4VO3Ld27acHX7Xq5jg7EYHsVzX70ZxXeUMcKR02gnhHjyEjApam3cSS3Io
jt3A7IzYa4tDVvQda3oyZ1OMsZulzDuYysORb6JkjWb6G7Nyf3732QRUES+ovd1R/IZyhen7LNUn
gSxNVQcjdK7xEWFMiINXgSBOTRxb7AAyA/idkTcXBOglPJrz2AlG1vD3gk//OnuX1gGRp+LySmTQ
sX48VuMe/B/Wv9RO6ubGt5dWOILb8GceJH4Rp/kE1cU2VwghJQ0xlTovKtx1Rd6u9+bpJfWHF62y
a/96XwMm3bZmrEC/R4AORlM+PA3gNhFZnSSQ3BOpmlNgPju4jL2KHVjRiScWkIr7c9GJOKEy0+0R
SglmrPtgLT1KHSh+RrNHQCbZoR2JGqJBkXO6amTVLGdclj0CSfCi7OwAxRZ+NZmuQ0T8awVqiQDS
fQt257Vw/bld98QnCZsgIiDUad+grTI4HOP0ZEEX7GMGrTlD0mfAK0fS3SAFGCKQthfiT45tkQCM
/F2YlQ/9t9YSD+S+k0YGV0yZfdAhzQzkKD7IXz1R99xhZAGlMbC/XeQs780PzZZhld64IHypyEZX
P5mfuX+KjIEpLkJ9Io//R3WSlyRRcjwzNrRYTynWnQwQ6VDxMVGeRnWIgWW/2r45KAfjkao9z/9S
rxlrS4UIZNuSawvHiQPX4j+10hW/MFI6meeGN2akVtMhlDMDQrUYS9RFaZ+7xerxwChNtmPN2XxI
cQXIjuftI6vtmO1Th0xXha8xj8fJN8zOfK0nVkS1k8HfOHzaTGSIZ299RsPhfc1QqfSE+Ux3jzLI
1HYW28oJSKIirT2XdHNVnmwEb3/S4bBsNFllx3mGHJdOOinlgoGLv5yWouQ3W2DGwy5ndGLWCbV8
7GnenAgOG0hQYxApv+QFYgDsTXBF9lDpo12xDyfiIP54bDG2rwOEPRbxckKCU8sIEqGDL7Nsdplt
wQrQeLkkCeUTTZAqQ21Z4bIT8hROfzVmVs20H8XEL7CA745dpGeJ2MYvMW2Ap+TLm6jL6XtgkELR
6O5BZtdygCpeHzL7OiFeuAoFCQ2HPo3/2U6iOMWST8WC/S5YKjQNd9RPsVY1q4JHdKL0YJlnzVlO
knq62Dj4G/BLCwfwoaM3KvU9FeAotyv2FudHGD8e4zkGikPJKdz/gR+5suxx2SEePQ54CEnywzoP
3PjGswtewgHy1604kneIoIMDgSobVbPcu444w5EjN0Q2lu3OPq9pYP6v9RoLAEY+xWYjWVs3zUhy
fgrD/Jou/XvkTW2Q9bV8Utc8Ew/GARJGte9zX4c2qXg6p3wIDLzpK8KAk09Xj5K086Zc28eW+vsV
9Yf7/1G79yClZevQOKAwEV5EnYPMprKgDL8WnotXy5FUYTK094rpOHGRSFiVxJHAWWJyHsXbFkE9
S3NCDUR7J4jbTLrpSXAYmGItufcbb31TOqEU4hXkkrj8SY5Wo8oBktqob6vYmF10sUK3nOBAIaUy
g2O7HsEgnUBvje+dCp9tVAwEnGHcb3PdlgsJ8tEDqRFDhrJ8XJquJnMZrmX8JbMC3SCnco3IMtP3
hcOExILYeqAS7Y9g5SK4q+/ak11SYn0UD6cQ1UsHN8mtgYDInbEHblcm2LPvjqCOgRRmbBxK6Z/j
OxpQEpDn5V+yprbgi57gh1Fn/uqBgBZ7My41iKQM5GNrByGjWJNRflZ2ljjUtL2+q4ojGk02jeJT
DLEulHK3Byr+Mrzie+QEDaNtCvFxM1Sfga2hrxESBdElJvUvD5UXOD4rkORcc47ZV9yCZ+a7QIDZ
xHFbTeByzb1nKsrO5yah9TIJxajpODzTPJbNc5RIYuyaF6ft8DkOe7w10kLaWhC4Ha4OkqsoYcwC
I0JfkMmJ7pC62U0QJyGiPSJ7har+PiQUA0u6OiC6LL9OdFlpk3awTHQLM671mjq8E7ldB2m9HK2a
Vm16zrQaZ4Bi+pG1YqFN9NZ4KW6nyyQlDk+z1anbHQdJuQpSqgmZl4UG5Q9S50lGbDjebQyKzQN+
4N2GA7Aqs86QL5k8hjZpGUIAuLEO8pwVng30VZvjWiR0cdHzvDaXE9JwNGByhrdeqKsg5h1rw3q+
bYw3BV6Q/tAjo5nTd2ctFufKnAip669Q7eA5M8qnDuy/M7Jw24fZl3zhvTeIsbCkgdU5ACcwbSZP
+L/6iV4OIyvE5KKRh5ndG55AknCZ6Jq2ogVTX7A8PWE1exkXC/+NJErRIM9vDB35685tcgFwg1vF
zn+47AKUgZvIbS6RIhhnKW0DugFquLyyzHgozgewgTBIKwEi0VRd+tGWXSq4FCIwBme3t94308/s
3Fmk6w3QOEdQqAuAKi5Vzt+12NwJoA3IyyT4jvPmAE64DuLyrQmeIhg6EvhLl0f6boc/W8klzz8L
rvUIv5Ijld4bPLqrLFbQRsADXliFzJakqvMVp7WdpIXnqlNUCbV0M9+mVaPmYFWJUlzCth/mgIaj
Laf3Lrvm8rP+NCoohCQLTpl408O4Y9NPsQzKzd7LHI5zamLKTM0wAPF6Kp1EyzaZzt8ZLzhwmos9
P48mldr3nnxIf1uT+ExSFYmrY9nbi91BKjZn0iW5un19C3uqB1e0wPEepAHWRqZ/s4vvNbCh5F/2
VwDbOccuUMDYwgPRxNl3fSXXi8YEftprSLCEDwmuBVfL4eP4SAUIKBidoa0CpiwKpBLtyIMBPQWi
YexretdBv6ZbQpxFxTHO+RZhuPyzy3pZswUP55llXghInGr1drwXgiTkVC40Yvb4z7HOxNrGY8P0
pJPK38nKn+hf2Lr/APp8TCJxo1ObqZgHpo2XjNGoZRBzvMRuVI6MAe69H6QcwcWPP47O9tLmMS5Q
6Z+yD6ih6vtdbVlLJ+o+ei0imgVd1eKw1qOKuq31UW+sS3/Z/CmwTOZzKcIvKScGo+RcrjlM9/qP
MAu/lTZIVc3JvoqmgsFADLPoVLFnwKxDDmAE1HVOnIhyH/2eGMfVvggz9bVa20Xr5/0ksHHhohUt
mIcTFCHUcV1OZY1l5XSqT+wgY6dPGdz3yK+UK26D0XqNMKAIJWym3L6Fy2TYGpIGJNErCLPu5FHR
SAQXbybp1YIWWELsTOzX3jio6+PKk4edZwPwSF1mVYQbITHv9z9D+YRnYSzaXYwMr/Cxtp5QzqYv
IZI/LKbDl4ywrJ3lGCS8Vobi10tm6q9OIKNrCbpNvctWb158qkhkmII/JpU+f1Rp9lEgWYT6q/3v
kolDkIZLqfhWf6EV6p0h1LXZPuQN9oVvwU0GluPfAAEDf4q0ReJOAT9hXisJ/7GXS96ujuytJHWY
5Ou1vCbKvVrK0xE+4/0Lgqs0TFWe7kvuAWyIfPuhtzo3rewA79gIRvL4QmO3TCA/23t8ei3s8Ohe
KHByzf/ivWWwf0SdS+HqgI2u77lG2HMDEX6a9sg6FWQtTY/L0vpw9swYOsvzHj4+Cd7emY/DjpGk
bRTMgQbjS07H64enFaM2Qh/93i/r/LP073VKedKpglXx/T500kMdzyzGf7HotKpdhFCYGTRJxgJ7
uqYuyq2jiYzdgggTDKC/dBMIxZryTtzoAqf2/0rqCX7aq209khjioZmjNXOyDYDBQLDaB+jOGuHC
kvOmP6l8IjqcM7ja1PoB2CbxTWYW1ASh+MWjHS1uM8DO1CXJ9Yd2BLmQwKDelYzA2+iJxrjECSuK
HmcKvwuNG9AmC2hHydECxR7b7LgmVvFDSwnbvPdI9D7ZKImfELQHGx9B6Xpdw3vAk2uLVd/T1es/
3fAg9yxaD2rH517FF4W/anX6dC/ErCYW/UonpMhslDjeHt/ko9/L/cTmWApoHMrlLlK2VZ8lJyYg
szlQDxIn/QLwJPqTLEasMlwBXk2l7th9oroAHkztmY0AwKRAa/y8Eo+Gu8sUdk5Z9h9bKkj5WKGV
F9h73hW+9zw73qjIFqWYQmG52jQ4Z+jPqejnosyOrpYdtP38QLMankZTVUqqbCnxwUMxqN2qXJNQ
ITVHbSlFX/ohMXcHIgcpWuscR+HyezIsq+h+M7vg0F4Wiveb1CeGBqH0C3T/qLtv591AuE7kxSQY
mCeiTVM+7Db1KCHJuLbHxA5AqMA3zc3BVt7FRS29/ErmttANYEGhmOFo4IIk+XVPby71fFbnISXE
BICEEBmBGs8nfHaJmkd6etv6EOkwsx34Hs/RHV+dW0KMDs3IFfpN1ew9rviQTABPC36R9ySdXxFy
q0FL+A7Gw066BxbuYfet63oQH7MQIovJ75zZLAX6+lHuJSkH1mDwp49jYeJSmSNqexBZJWxCg052
7pJiVTY6BYGF/ocxE9fjbPDrMso1r9pFy6SaDRiv4IWyORk2ZBqsj0d+Tlod7Thet5GEsdzM3ypc
YVHUgJvSGutoQsNHUmb9ShN6jRc0x4OaZ6iNMLWJ+FoUpVnl2iPxKMQZZakMWSSQtpADBo9FoSBV
OTvr2EvCzTxg9m6MliMcRMGHLKjqOJMdLqHC+pe7AoX+Bp8hVO3T9FN/lIiJVFlG5ndZXsz0ZjJI
h9+AgutqDwyMbynehOhHXYtzI2X2nbsZVhV7rIhHG8ntodFAKggN96biruy5ZXF5CHnRO9omBued
pG7kFEljtrBUIo7x/KhH7sJZ0jeviUmuI9fRY++b7lGvq7boTfsLaJEuHSsECu6rdWfpCguDXDNB
e9i8LI0jhxZcNlk5wiZQDZP8rOZRo2ePxPVyTdVQqRnTfteyjcF85htiGKhguOyLz+rY4tu+AlKQ
freFCDrIa42LHv93SsiVipFlzc7iC6ovT1vLpzEaU1Z7XAcmFAgFokRxaB1S38Wpk2tcgINLneNG
LrXoEcI5BNHHmkHa7yWmW6D2hgBuRqn1Qlya/FRwg8+nBJzmqaR6eD9sYxDOG5dwfNWVQlz1FUWl
aQa0Up4tG+DTrpJ6Q172/RLPBVmPHyyJmfPjRz+X9bRVvf5tVctq7o/+cFspkTlRSF+Q3twg1SNp
W345OZBWZkzdO13f6M254PIPLjZv0BSL4TI7KrM9COte0V8N+JlV8fcWq+LLCLnCVvohpCjF1WYq
SWdI54tYfNo4EIkU7w/uJKzfmbIVq3N9xIYehRl596SC2kP8xfILBZD7Me/V4eKQtLDs5mGC2e1A
59zzm8Fa6l3jziAxZTO2KttHMEmgl6c72hTlkGQ8dmrB5VIT+PKB78jDkkpH7euWULz2gl6JNZ9l
7Pr+WfXsYYIR7In2UbsqUo7WkLX6oJ2Lmv1JyZW+CkFzK0E5eZ739+Dp2rqk5Rj7EUP0YSoM5kID
cL4JU068XuZejeORdCeZP5apy46PYEX2XyJDsOmBQZUTIAqcP5RVloIEO+FBi3MPQ5eEjncgPfKw
7/JNjddIx3K+ncaHMnX89pxqT0PwFMgoOG8Hx+sqYu3Kd4A9IMeg/urUieTKUFVOQgAL+YnHaExg
goH0DovBpglZr+xMzHY/y1/F4JKVSFa/j1ndITS3FnlsJ0zBbhQ2cqqEcOOJy4k2dCXvxNVre2NT
1bmyWMrrlw2X7wiQEEjsSaJjH6BKBz82HWt+lGcSYDX9ZUZkOjF6fF0oTBUIyBu695K50MAvxylV
C8ryWknB2K8fTzgks5qdyc7upgu302Z6O+jpozdYVvRUnNbEOhzM6awlbn1U6ivMHKVohC3eYpd8
lRUbtqGidH/x7UXpKrmX4zPV2nnvdCzIhuHTulbRb3S4p9xepJr9kuNqg+cCXDYAocK66MHPxSFU
Y0B8CP7AXVPTG48KqIJou6p9S3J7SmHffEknYdIR+ag3BTnL/D4ue5D2126XBtBqKssKtzw9DBX1
lwt/OqUCN05VjQEYQaQNO+x3UxGk9K4qwqwHHhbSmG+rRDvNSUmNM+EJM7Hd9GIo30TRUu+XwfHn
E5uJMqgeeN28Hg0KW4y/a9wFKXOHiw/w0A5Nf+nzVT/pitPyZOxgnilNLYSr+qxaOCwJmVnRBjri
0maAeD/nauvLRYwVcaXPQSUCWdLnxfzjlW03rBDAae3hKFk6Ji+ULfIQRWr2aY5xVf0+yGSoy7LA
zsDhc/K3HoX+Y5o2BdHV8v5smVaBSUk57NkqD1GaHaOXSU9Xpzi+WpTQptF3f1pAGUe2U6IfC9oP
ziYwV9zlpt1snE+cl9weri/fl2x2VS8W4rWgqGLkNG7/O+bDsKT7UtbhizWmOABjVYuODOdDQJas
O0ZMuvedLbHXUOzYLXeFfDTTS3GzjzLQpZqwp3T92/KoTO4WBoS/alrwzVGf8xgi7IaiplCMv2vE
D67PBPg2OhQ6TqdgHJxCeTVzwnPPuhmeZwYQeOBMXgVdxvcRV5IR2k9mONMdZN7N+5h0gnDSLgfW
uSdqLuzXPocRlBAPHzL1/krxR+659I27AiZSRma5c0x23mvFMKxJJSJv+hcq1rc++KUMEo/zdAjM
c65QCG2IsDMgC75X6lBwmk8AO2hX8/ELb9q79gkd5OYlg0k86FVMu5NFe77EPpxEALxz1JdNuims
4Udq5Ntel0mi/PahYsLV0mdqSErqMU4GCbl4edPt6cnsEc8nFf9MJfm/n0Esan8pZfPj82n1Y23R
sJL3um3jXg5EAvHKi6BPEwX8hn+Gm4apsXx4DVgIhiCf7yaJrNDE4TOb6ARyHLQlCIzPtfjVh1U6
BmWKWWX/rRqHbVxhl0Z8xPwDPcbcWF9xmKTR2OfasusjCOp7oavDsHfSK+xUxeEFjkNnXBn5urVn
+ZkRu8EbMofdOBL0bmFXBULNsev3wXJPLUYyeHwkEdGgGwdPG/1l1MHbDqzq12EWxU0q+JL0ArxR
cqOmPs2B5e+0W/l6mnO+9UOQpeswe0bRB1CpZr4Ji4hvIDao5MqfwODTDHuzclAKyQ+WhT3cch6R
WKRp7d/UneHXtct2Y3KqsRrEKzlRp9/uedcmdJfSefVWBiHqFHPTbGUBHU8ZuUGBMpLvVHi4JV1s
rAFuhRz0PNF4LzGnHiDRoZu3K4sZ68qwggEFK4p9jNE9M/fRUqk/zX0ezb+ITv/nBDWkJvjfmHtH
gnrPDuoPZXhTQcHW4ipHypj2vVojMP4OO01Tnfq3zLdVERfJLuDi1qDn+KQsj9I4GfnznCROuxR3
G2QOrf9nw5XN0oxIijdadSTd7PVCghX3VqqxbjjOx7v5xZefG3pRMj9H8QlcsUlsMXlpbn0p8Qfb
th71RP/pgKzj2ZXfQw8WgHt7xUIAWe2WMdLYeTysvVF9TMIP9YpnxFh3bI0bK3+TtLGyemUm5301
f4WrnKgY2QjHp+6IBZV1mFWVsUd0OwVLMth+z/phfSstcG7XNwS+iE3915xQG6lguvZqULpTywua
+ZJ4gcaB6dNgXcDJtykwB7Hf6RsNM20lKw1eoZ9ev90s7MxACYyn7ELig9RLcDwFDwR2xwHL+7B9
XmtyngpCoIm+NY3UXUG31HM+fe7kSI7l+20DHUYhDGqIxp4NvrM5tjpduzPBRkODXcHyn/HCeRLA
hfkAWU5+Uf6+afJBEd3zBJiK66syGC1OOu75KhdPPDcofianHerd64fKPHX6Bm1YD8AQMs4mYKIo
Vwoclt3cKcr6eWK0xQssZ1Yod8niBsOoF4HXxqTto3LN/OZJlImLnlJPbvrkm2EmX/0Gjw7gTFA3
zYQt8rzEpSrpg6He+QuKkc1mnv3uErL8bK7/Q9RLenoHCEsov8vep3lGpjafy9EFlJrdHDJzNJHZ
2xR/NXghOfkoEUhAA42FUCbaMsmlGTMx62cnrcjbkrgnMDwLwmwBE+wl9zEvAgoHrBTKDhnfuImq
KSRS5UGiJc0SsAYEoyE17rFUA35VgzaRJLmxQvaiMIi4v4K/gzabvSVhHuX7VqUCcZZ5G7Y5j67P
eZeuO55IXUZJgdGHOi4NtbYFkAIUQFBGKrdJUGq2qpO6y2NPPu5OPzQlF6BIfv8gEJbovcMJ6Inh
KfQO0IsV4VTMRR/KvuhoYnvqqSK/RrWEx4eO+pk00QHFqXKTB8gq1HSy+BzXrYwUoAi9doXNn3Yz
9n3bV4vH2DNcc130bFYMQeaNuXk16ND8TmCopKSlxj4qOWHuVJQhkUIwF5nv94CrKx10H48Gi/Rv
fbo3X68IlVsJ+WItFDdtUKP8BxodiAaMGCiCIkySzw1KiyE4LiXRLy/B289HDlSWKMQ2jdAjX4Yt
esgEeErVd6rHjGNzzeSs4pB+B/+2ahhMr8vF9uQPwItF2Tix6dzpOy16zMi0txxxWJVHBR/Wbi+e
rmfE7rxtTHx8GkwOvgwG0DnjLJ+dg0iuUbBFJh4HRcfIcdOQePcLE/DsQLy8ktPwo6wGkeJNur0s
DK8YhHkARa0gPUtw/xstR8QxRuauMo/d9D9r0YTtvWFsfYBVh8/dEyY3ILmQGTdjq8Bol6bNQi9f
Zy1S1b1ELxlBy57PheS+WfYlsJyaDTzTV2kxPKKoDvswh/PtjfeL4KfLlrSuMOPwsEAn6gCaUqIN
m1B7ZtQKnW+xOmnjKzdM0VNylu73WRjKPhLJ/6ejWjwa3aq8HeJm8FiNvV0gLIEa++yCRzx8JiZ6
aZbxXE/K+JHJv2XYHz9fMefkUaNYwd9CrE3MZ4+VHpQ35T2SWoOcsyhXELAxn7BouKzPejfciVTF
5dhm/KvGk30PwzMHyYuu1s7Br/JRK+8N/S54I7v7dWao2VmvXDxZOgKQmt7L4d7VkjlYUtj3Evp6
RzZeVivzdtLlQaXpHRqyZD+teIZVbRq9hb7k5BikVwN7pFvwoFkNpYKZRVyg6kJjQmFFgRbjYirI
iZg3oePaImR/i/r+uagHbzAu6stok0NXiZweNydt7JuTw2lRqNhVzWavNGcQP5zRgyoq3rwumvHA
x1OIC269woaHagw/9ReZu/DzZE4pzh7jHApohX84SqnHN5SV5WHsdQR66ftQ49J5n2eMKSit2V3K
cX5SLIyg6ubbb/A1P0n6M+vEafR6l5urlIAzDsY/vRlWM7BZMcpIC8uNT3LSSu/r2BOfI7tIz+Z+
MfQ0eXg3nILGdCpQzSS4aCM0kCrEAxyaKl5419gMX1XwKGpZnqXbeK4LnG8n5NpzGec0OOwliNLO
3uPMz7x9UBrWRwEtulNwQAGenR95jKIWFgd4sVE5E6ulnLtNDhUbA5WhT1ZOoyAgCuJ2zALNeCxj
sn5mU+xWCVVlA6J7ZZKFRqwEXOA2Cjp51E/mBj2cS+DhraVr45Gr0anOHVWE/muF9QFLRRJYgRl9
yfVm8xeddVCv6jG8PhN1EHv8dsPzy+qMYmTh326A/QPd31oeWPELq7SCrqeLMwrKUFTsNvclAS69
77cuZSITskYK39viveKLxDbbLp5aMBvyG6i3u6I5XEnN2+5FyLQ7ACOzDvDeXHwoublOxJUJxVig
98hSwJ/HdnmEpzcJGJVFY11LxYR941/rR+3xqvtr7UbPEktRiJfdtAtVtPzIYncKW7t07/OUY5PZ
xhjUVR3ZPV/jAqUsXh1wMZOdom5Xp6UAQJWtP17sWhjQWiLGJT6s4DvhhTZ1hPFxdNLH1vRjje5g
zARL+My4t/c7fi4gZnZMn5FPdCsbn8LBEvKC9gvTvwgZdMsi12h+t0K41t4d6DS+h++NUE6rK/bE
yLnnxr352UdsStVkUcprKsDABHEK63b3bfkKD58+Z5Q2Q/NuAVmD4mfQdygD/pot0ym1JsLD7ZqM
Zb8Lbfgrc1v7ebRceM35HnAScWqI3D6o870kgvKzU4Wre+vAnS43o2h2GDn1PieQAPuujBNKyDng
zCK8lcXMgzK29ALh35xmuqoEJYxp5w4nYkTEwTK/+UtK3AEEC92G9Z3fc978xpSOp/HsZL5JHOAJ
K2mGofUSTkDPiuFmMP/g6qHRKcaeMDNKCTZUQPVxebFLNbG63u0noKEQy81OyrqyW/7/4vxu+7p0
+1rvDUSW4KfQTNUX2gOpLiOZMYMrT0bk20BHzcBwt2q0ow1mhmQXLj4Ejw2r48QxsIE9NKoKST//
QWr91Hjy35BXWuu6DI8gVBUy+7qgFBHp9vnCyrXTMGsCQ+h7YYeEpGb7z+M3Gh73FKQNC8gerXi/
2JKebNKMDzfyBq+RfKCBuAe5q9XJiK9Ev/b0K16y0va416Yhx8a9a0NztQvHWE9IcOFGpUEUoC5x
52Mxmj3z0h4ZIO3MZRfB1EzeI1y9iFXmAHxH4yqplHOKGrnqEqPqCR4yx1goeIjBizqlj27iBYLn
iITwXD3qmcvfe/F2K7LpSnz6hXXnk6S3B2QJNWNc/rWSY/B+fH6CobJXDSpCBlgkaN1h/ERIl10z
Wt8LLCgfoFhhiPHRwGJ+sppd3QfrVHZb8ElVxYu2lpiWydafnzsH6stVEeSQqxuIJqAbevZIDfIW
WMKVqf9jSCaC045lpqvxs88FGU9zJ7ys0csLX3riCvRkd3W+cI/zlHbsQsHfbeSOfUiYLDly7e8b
2/5YZOG64Ez9P8f6iI7oW+cPFiYbob3e9RV3R7HDXQUtAFm8ZY3MCGybCfLwnzdqxR92gcJztXSK
zWK6Kg5Ts5yq91deNbKjcOtzLxt56pVTeTmaLrYH4uzM0fjrJba8lREX+b/sB32Gz1eCnpsdS1Bq
2kJKaUpbJtDVfEY0YGgk5IJ5ID3Y/eABF9wOOOUlBF1eufojdFw+sJMGbu6bpGJl+YusDrCXyuoc
LFZxVUV7b1fFDLPUfAJFSpzXmZ+UrlefAeFnsyxQVFoyPGWh50ELR2gNUJ7dWJD8Oo44BYfGEod3
5qckJDBU85YFii9Yb1pCVMXuTBAd8Kpojj5WbC1esT3cujU/kVzuS79w4PTngX/8UKsQd+aaxmsQ
8mgXUjoNBFVt2Tj5xkRYaJQCO/oqHEFF/qnOSo43IuxidIx41AMiNOokFnJTyPYXukOlFTR4AQ4q
A/0wHRswEepgY98ORBqhUC8qMBNvpddyrp1xGHKS99Snl3xve5eh6Wl8eGLG0oREKcB3wUOxHOvD
x5Os4Y1QivVPpEnPFbXqTXFwMDHJZmCEiV3GRnioLfrz/Wdk3y1Lrddo9A8/r8afyxM1oFCKuNI6
kCGhk8S5+OE26nqDeKkb0KI/bp1EJlQhm4yZ7ZUFbvuE4b/QkMYkIgVnfTu/JOaOvp2Rm2S177an
XfXWq8F49aCqswtGARmTSJxd4efuNZfU/UzDhD3J6aINHOwKmmPefCt7zUT3qGqLLB0e2MQVIgoB
MF2PD+cTpqbJC+L91kXZkN3rSEfTIWuKoffKWu0nPgyy+H8sZVyeP1GwkRNWyQwoL1NleC64ayvn
CajeiHlT8TstIwORvhqTUXgJGwPp1zcNz+SNFGV5AeP442aclLsxk0OD2hBy7D2aEkQheTUyFopF
FXi0teJbablgU4bKbgs6FtYRMtrU3TMdonTvnEIUsFTtorS1xXyrXIm8x/CKJYe78mDFTRK5ErAk
ZmK0mVfFMWaohiJVrK+YaFJFSO9KwWDg8MNgIAyzoldf4M0r+iAgtypnspTu/gx0GpX8MKkv3MYf
dTpYS2OoK+HgFv4cTrhRoWx1+EWOpKTxZUxFXgKqppbLU4MTZRaUvZteR2nbVA5MuK2g4c3uEVfB
fp9d1dsdUSYQfLF3dg8t0nPPQCr8NUNzoHAh8NeWX1R+d0qh+qymWmPZ7ZuQP2jmxkSkCgvYzN9V
hoMDG1/irwHpiXDn3joyXyh9As/SP4muxyTivUOtVYva01v/NP8KLmxuyEfmLkkbh0fRcn68kh9M
jL7L3Pdn2uAYlOWrPAiqqvRN2b9nTzI+0WRmBEx/lAbd1JaJtQ9XaVNzCeqahZZOt3PYIpfYLUnQ
zJqH67UdU9PsqkiGrhXpXBi1s7XaMqu6n4Zw1hpbDYc0b6AW0xelZopoWQsgXSrOkZmqKXrB0XN4
f9BpunkudNrGuJhZdwGkDBDw2OG72hfy7yoLmfHSV6URnc+qRtSdaqLepEOt3eETNywrOKC8F4Gd
bc+YbC87TZlQJZN50mKMMZis7g4XFrt1IUZcbONkkyC/fv/5bwNd2Kj3VQNrcoSzPSQOMp2g0KcF
69xrcCv5eu6OukOY6cH8jLeUBKModjfMlZz3z4cju+nb6eSAbi5OuXOt5HhAdzSKmjVOFpf2LOT6
AVTxUhJfwKQDEU9wlKsOh6yBocwJuwR9+zKqrKMlsVz9jN6VRlqFlOtKwlijhCkIYv28HHsOftkc
4ke8+bJ3vcYUxNaOwuWsgZfyTRlygmYpfpFFIbiLDwM3CnS+rbfWs0irIWmk+4y65i9M5aa3QgUK
xQVrOeHPrxjDW5jYE1E9pAHdWiUSAEwnvrtlwh3SAF9+GL1/b4hT1GTnBYOM96Fuj5pskzDMmvRM
5H3/LVAKtRH8aNBaHinyzCXlvamGKGzmUtArz+EpYn+gPAEu6Ac/LFUCQw2e0j96uoqFPXtNXFhA
IFiQ3v4wgrb/xgkSOGrKV7kwy8tPrs//0P61mQXg9vWvTN8Ozf43qK5HdCbnR1VV09OJIMQpsjis
tARao2CzevaOlOGFxTcbZw3UqwId7fF3VzJQEtq58hVdK4B3GikKolz6VoOMPcTcP75vi8CpbRnt
wHfqLtXRhKjB9EV7wQOrmRVze354LJWdH64XdW26r3Qf37B9E74i+KdWF7ofi57zmPVBsCN/Dk9t
PZD4WTe9tnvWm/Hnk1clgB8+xCdLaYGPk73xLg+r/IDKSoAwgWO7vNOkTm9QsJMFEtmuVnS7Npi0
/TXMNkpy02GGkKmT/D0VSWro38aZK+qImsfM2uWk71vgRcCL3IPFrIij9JHeoA7yqzth+VUYCul5
6yPBSwT0WY3TT69XrriDKHSEQ55n7jVARrfdX1hAASnwMGGAR02bBivsuKSgi02QfRcRF8vHcXwV
tiykucQ9EsUIZO6e+R4dHj9zWk+mMud6cWI6q1XyzqRiZTNixNFwRvPjR/EHdFKkqTn6UNO5ceMS
om8iUG+2/NqGVkj72MXJ3FL4Jp2nF/4/0VB6PgxE6OucMT2KeygugnMvh6TaRuVdWwdIXiM4E5/n
yblILSKCcy4Ej5qSk7DdH/ucp05rWhMreIHZ9Gxp2fxSzZYEf/7v5swo2Nj5KgyENB7wpRKFNoj2
orehRGEJfVqjVV1xSYLX39KAWkMN6Z0ZSlm//RKHtruDeZ1CGMEQE0gd34lHhfec3pVy0vijyV7R
60G4HLUar2jnRyluWKKFT4ZkTKq+kIKr3ntEHDt7X0i8RDEoOZQMXXGj9fBWAzselgd0K+NE1FS4
tyadOA8XdIZ7B97AdCSPfTy1GN+PV25pEU+6p9s1DiT79hDPbsFB+7Cb2FTmcHETW49cdqFZo32l
5D5dk18DnqKqpX6Fm27kr49gU/7NynAQ/dsErJypM4s3D2XO1vQsF6IzEc6k9jP0iDy0qdPV9DmC
fJzJR77JFBRR3ZV7cBAXKiMdbRF3ve93eFll37mcd0X4AldK1Cj9UL0ZuryxwB+EOBxDxsLmLWaz
EGKgK2LTdwr6HhpqRgd67f0DQo96twv233IO+uqsHLz+ONHJpPmb4hKDTdOuzB/Zd5sLOvqXLkLR
ID880bLY+UwnQ7lCB6fjljmQJ4FAEgdMeZ2WjUpjMSHLApXcp7DR+0ME74Q/vNMQCXqY0NGPEn6e
eIcKqiC12ZwhAfmDDE968yGDBGLi86pFOp/rtALyZbdvnP4e+pOm7O1Ij6beiY+ctAs8NOfJ6ocG
EDmbSA9aKqam64EZqgUg8g4bTXGRPOuF8IpYOYpYuZftm61tQit6w/w9xYGrm7g9X5ILaiPGsigu
MBHCZ7II62kr3A3vl6qbgQdC3jICLfa8QdDaNkt+QDcn0gD8nuor7mdy9zQxlk879heCTrPp5Gud
wAKLVSyZXT7PV+AY1uhYsdgdF6KBfZonj0sy1pgEpHRCSQENVckh5bNoJKQVQ5oB017NMHMsqRGX
SQYiKlqh9E4Sq74KwNKK0WeWe1L4jOG4JFRaCAPfq90jURNHkMPcHhrmlEzNjlW4HuWaPJCt1xvQ
tkwcpsUc4mq3StdWZCyhL/nTJeJeAjFY7+lW5zFEwSmbdORsxjEOr/tkMKhXogWRunnarlRB5koR
i1vOujojod99q9S3yzXFW6ccC01eCc3CGh3dV2+sUv8cgujpufQOrdqaD2Ij7YFe9P5N99B8ksy6
E8KGJixR+3f+e/kFOiJxPkdMvJrKXXttacXcFDVwsi4vT+q/LhrRmIxds3/j72Zx0NgU3h576rYl
GZXEjLMn2KyDVvahCpDjKFQrSyEJMZh6usTT39vdtjoZS6VirS3XAT9IAZHmFkjSeUozAGtEZQDA
jBHsiP8PtAPAq+b2FWLbC9AQ0CbUd220w/zVUvcsNEcBshx+ss1++FVF3zBqr9ax8cNaReDoZ7Zp
aBuw9JrjsNN1lER5CzemGydMxoy+8AP5gVOk0jjA0wP/3IDr0/WkV4boSIKssak3ZDb9nkBkzlJd
3Xsn13UlpnDR9u7r0twEHZhvsoGc0LpewtyCqWSHJYtfsUBvlTIXHrtSz4Eqr7af3j71SJYjfKu6
pZEywyna99O54DZPChNgpmyt8jmMzXalqeYsU2Un5yI8W+0hKCr5fN8JOQHoAXMHGq0/aSmNT8D3
mg9gNBfr56L1K2sPU8hwXR/V7z00orN8FWG4udAKuVw33o/1EFcpOADRLJdbFvWMnOSs5zw5pQOH
5/Bq3GofcJTWfHB3gADSuQq9fY2OCg2XVei9hVD5FthivEBDljDIxKeFFy0sRKaFGYWC7Ptdtwk5
sLESQ2Pn4pT738iulpdnp5kVyEBzFtdm2epitRltXe+zpszu837unVVooO++67Nl1f5V8deXw+mZ
F/pelyGqmUYlABmsGXm6smNemF29dLfWUkiRunek8bc+Y9uUaBYvxdg3fRVQjGDPNgixLhhLOGbu
d+8lXW4Jb7oqVDvcZN5Ym5U67k7ocyWVmhhPQQZqOwKPMJ4sBmet5gxr90WlnKrSJcEQmwwVph09
yhvMDnioxPBVGdRaikNObz0bnpDKZpde66ktWaBaPmUc+7D6VUMap2+gf/GtmiEXfplthUbubZMS
C+aR/Zfbt8iRWWBrqwAnDdu3GwdqxXrunX8Hsw59a2t1a0qoGWTL9nh2hyU8Sv50U10HDcN1SFmw
4joSJiYaNVbSH1r6cnzYBzU2h2M6sVI70WxvLebLC7bZ8yQHIjNZLvJLtubYmDPOrxUK0AZsOdT1
t2PJypwva32yfTy6xpG8po477tMrQbQxYeA/XPinWMvjlHq+2oX6iCgc0YXSkEldS/jpkUZIl631
RznF/ST4Ty3NN+kSpNhDsYAPWz0ppS+ORt4U/Dozlf0pOdavTKnw3pm2KtBhyMPJPNwF9ROXIe2x
DLkWPUVk+HZhcq11dx6szzN/3A3Ea7jwUqgyZfMdwP8M3e5IsGyNdps1PPFnN4QQLzlnIxuQKuLd
QkXvKkD0fIBsu3JWdUcWHefbfz+sU+Bnszr2sV+c5rt2KRrs6QhLMWr41ADvIb3ZI9LJhwgPwRqm
JUqaAylA5XDCfEy8G1RCxiofavUXqbjMkeOgiclLgf8d23qJtUhlrD1HOVkYG5unRy5zaMGZhmRL
lD+xXFdsojOWStdUhAJhlqejG/ezlgere/Cb1+DE8Pnrhq6cwK1aB496POSpd74CgMC1DT7UMCn9
g3dBb0qxNPyz9LNpgjrOYtdeXX7Vb96tadh9wBeA9lfzUIK0QhpY8OtxbK+/Pc3dldR7TCCfd5tB
grd7S9wut2LQ8ja18JsPFOMEppGAzSdc7qk10xxwNs18BbptWrsUzOH1/awjewoJazRPJjoiI1yV
DoHdwCgp1+g4frRAsKyNEJldEpEqRmNlwfNTo+iqzeSghteuKXp1PVjNSfPDfsKN6UUAnob/gfG9
VEmwVLk1LWsXonHejPtaqe6hurLz49BAHqGXXWAgagCVEM2jHnzUsH+pd/R0Sblry5vACrQSuZRr
KEXVYtLqMTO2OSwETkrwlCelB1ZUxIYEXMSPcucLpXU4N3frhGToVpaHv+9k4OpAh2bTu8LeIaej
iE9Ic49oLW+suLOziYDYT0brjlvNXPyistXioMf9URClbhT1O7hFloth01jyB/V1OkASe9d+bLKt
2c1LGd/j2bvM5yz6knGyXPAwxrCsajMZW/vFEbY5iZApSa11Yb3BoS4pTaQM4G+xD/CdVGjf6vUY
6+3rhy5SzeKXyjbgNDC2TjXP528GI8g5QLhJX6Wz+EWqzMsDLJdCwJh5S3Z692zbvqVvSZrBwF9F
eknt9k9brmez2RbacjheJPEOgAu5S7MkI1Uc0eCXgVBhSLRqpjYWmQyHMrUJveeVSMQ+OhjekIHC
Pl0xTEYyPSlpMmHfSk4R5W+wlsYEQkOod/ki3/CkMX+k9KTguagpmmS39pscEwL0PvJUcKkK4Eni
p54NqVUTujl2Ik0v+B0SthAbPg/hPkYl3SBkLsnJU5thCeldz4ZWnuCYY9TYkaiLUstRbQBuq9cn
6EQcRtxgVCg8s6ODWKeCQQj4kuG3BPyA9R7WZCmij92RPvSgEOsxdz+3HsAOMkS+FD2flh7nQXqs
dREP1sKOl64Q89iNA4J3AX2db6RA/FEr8WJSUDGIKWTl1zFbpbs40+1C3YeAEH3qZkwaH2ICXSpJ
CZssp0GtBh/1yxryjqxiwwAxm2ESWAMCl/WW8LzLdR1uPHDt6M2w+iquWD5tLsSfa1JaG5S5NZkl
mTjVMoVR7CpCmuC555CU2dfl/QRWswgYGJOpLg9ZpjT4l72D9VHOvUYgM+3zVOA897w8odk30N42
qhx5mVeTzX5C0pElfsEYX4W58xgXVHkZolVtwib3ELnjj21uKA+c3T1Pwqrg7a1xZEgSSqnVec8J
a4X8lqXITtTUQevcf5JgatPyyiXjFhcuSoqdFXz3ftZKybbmI+or91GIbll/YFAPmBnjdz9RQA/+
9pXUNPqEHzhKRq4Kzx+Qk0zQqm51N73JLqOXT5/vEpHb/VvTRB+Au6JmN13LjrvcZbMgCtptj/yu
Xx+97A7DOXKc+8zf0NmFWDCSAQl/MQ1ayju7T5dZMFasuc16GTinAHp1eT5Slhal/ZEEqF4uq9Uo
j1d6nL31Ym8ish5KVr/x6GMw9bEfUfYwMlHPj/pBMXz6BJNq13ZeFCIqpJib9+fDq9/OEj5ExCkg
ZFzmqRvN6kKeVOKUpg23XfhYzKEgaFI40yesg9DIuVmOth3/+nKOXsCyF6LWeL5CU7SFoH+dAsho
JmNCsL3sYoVjDn1EQrkZxXfZeowW/lJ2dEsUYFoC4fQf+Iloka0gKLVzCEL6e0/sIzJm3LBqUwwU
eThmJm+K9JSTj2ZKCR9NoPlMLNYMMb6qy2uIjUO/kq1XomJyUb/EMTjmQzUibJhzse4QN1NHf9ZP
ZWFboDTkvX1m7gRPCpEZKlWJE+vioKvzO7ywSW3/FmndC5beREH9JOm1Yckv55p3HqSx++PaKo48
qIRfXNnn6x8DBvzpvonewVH7Q/nGnrf5UxA7OSGR6zrFxdPtCs82E5/zS8LqXZHNUlZ1/Egmw8mV
bEVpTei3Ic9xu0iNIPbsNBZVf1tmPn3Z6xcS4e6XqL0ZxHw00Zzg7HhBXgsWSa6abIH9eYVcC0mY
1fvddarA/IDiDFapkP43zyMk7CUCHVTd1Ytq5ZtFEgADrbWW4yMVInUZTiSCI5v/lmMBQWtWbnbH
q6Fit27Iazt9Mm+0sQ8mxIwLYs5qnFbaltQYI4OHz/MGGexaaZqfxVB0o/lm1zzrXH4RROTH16R/
U3zNdxhOmLkA4KCEY49D0pPcgObwX78Q1hDgrZccFOhd6aOKf7u2onDAtUozjdJCPjnRxmn8rY4o
EWZNjKb/vQBILVZ1oe7OtEBcUmymH4BPO1N9Iis/YWHqLYm09BI+8/tRpNdzgYd6F0MCzVThxPfj
kRbkTepBzD12KsE4Xt9fIw4xjk5wcVCJJZbJRG8MpAUWyS6Aoev5F4/OKeX368pv568YaBW7KDPR
3cjhThJD+a/IqBzzzuPIuSzWDjMQNtIHA6Y1sHewGhUz/4tBPSrRFl3aYBs39QSYWVyDL39OfXNl
Rqd/h2VUDqhhjcWYpU6p0ylsS/rgdkmLb0eEP/u1vsNiL3ox8kfuMLhhbM7TTsu0ydkYg5nsrEPb
BvSlDFNxBthOYjqpBBqExQaMRis5c2NDJnHmYrG1TsR4a5eKYtCFtoXIWCd/SHFrvAzgGGWms2w+
kDLG5wQv9yO922FxkwjMLyB7+MLDcXmfExD3PM2rvTgLfn3E+Ua8NtWdF4nX0SWvPrRTYqwws2FX
R5Swd8tMKrjxa6yjtK+dq8eIniFcdlWdq0YItfh0dGsxf2KNFZ9ppRV3ZNrq5ipDGUS7cLeEHgPl
kJPd9jkBaTAL9iogdZYqOC8PN0RhBs6b3OlAZbviK53kKLoAPE7OuggQnhE5zM5diN9jJs1RSVNe
Mp8EPQilejD666ne+MNtu0Y/Lqwi5s2iiC8wElP72vJqPqhPxo10gO3ZYFEOSa8Ti/4iL4j9LjUe
CZR7CufkL81OOiHWEp3vPwWy+9XyAi8B3oxPdeOW7p1rFzeUB5Q0yTYCvPu1Xw6WVB8jY1l+PVLa
8Etc+3lExbUuGSEUReq+Oy6y6wWU+AOyQOuY8Kf9HuPX+vn8mSyLdww+jfXOTGT7RxTsYiCjBuFw
JNw2nIlEPmn7gcAR2XNafNvfdPnwDGEY9rpyHRBZP12AbDfOZOjVx/GZEmTBJnga20L9ebtxwyPX
3wUgByzI+fEeFRGPud/cL9lM5sIyVglvomYGLOuEpKcCr82kxhhHFcaDKpiwPCjVq/kPcY9uuan2
glHNaWZGVCeRdlOrbvr7EhomXd3Zo/Fa1M6o8Eq7rM2oCZqDaa4b3rIrJiGQBLBnmWem0GKJoLfq
tTIHlSLUXn6HfQzCDX2h0OBrvsZoo0iLW+NvSbSCpf5odn53ZxcpyVwk86UgLyg4HLM4WXgCN768
64lf5kwjCYXnzcfdxOpIgc9pB5Tk/N0z8C/b/grJWzmVUbNiTj7WaxgAlHFZwiC/41YODkWuQF99
ZAPI+yg/AgQYnvkhbW5FLP3nDex3UVeAucpHQUCibNdFA3nFgRo8/NFy5tBuMm3dVvBUFUGxJ0X4
XsLtLWuxxzqe1V/EQY7Jy5VDx4jowNTSqgDqgtw30HXQFcGJihD4GgqxQg7/RHgSOhgKhf8wQ+RL
FIOOrQhaW4h940m8Q8BYWeLDQpIqotm3+VyvHIRSQKd4GAe7GPUWl/o7ALX+ZX7RfTeWso9LJAlU
k2CAGuT+rFr9Bs3TMNIvVCBPc9aT0sLdr5IbH5CAMXri03AJj5dOhnDIMGTwKPdjSiwOi9G9annl
W6vm6ewfcQ5FeOOZNmzE80ZQ2h1T13LzNr7OVmQxQ/1yX5O4q+9p2Jy8cCjwrOz1k9mOYWpR3JAw
hsfDVWqxQ/Zlwrhc4wS8uC4Y8CQbiKxAqts1eP809iuc4M9cHXXMgDdartvNI/wzy6EbBmPPXRkA
IsaLuBaj7gJv70lzOkQqjneWeRjZHDmWEyOlb8wN6rkRivTxcq3i4vUrBwOpuCLymFTIn56ABlwP
WUnIRyQfXJSqDktDZxejx5uuWC7Iou/4LBfG2+YeBU6U1e85uv6+CUiAcdEdztdgHtAntzXC06kl
7X2f48bTPlE8fFsGgrBKirhZSbkKhePyAJ6cTs2bFEcRejS3p9epDF2XGtCtxakRTI0YhulXt+Yw
XdmqYqbkl1p+CYwsxfsuwekNt59yDkLMpC8aBww5PhaovyYmVWOaXi2BArsfqhOpWSEkEHuTOEZ+
zO0BjumDTHvHpTnxibhamz7W8Z3oDY9FlUHXUp7N3l0pRBw8Nbb4112gH/5HUji08PDLTx3LeRH0
docgtkSCUJtgWY31lnXAdY3KZlYWiS0w2rMy67Ph2BlFd900ZNzhvETAUisMw6OCGMJBYElE7dzq
KSwDat287RT1xyXqjSKqt94vXalnFHzrWzLiP34ut3Fbgrf0fCoD4Xoifq49eb60y82zVpOL2K1P
fcM8XNSoupZYHBqmJBO5RHuHx5U9SrwQW7qAjOu+v0UQX8dD82vuGFT7esiHzkGk/q4OVf49Ia0J
jcAZ8Fl/t1bUrGzWsPkC62IAtTqsesuUWO+Qqtau7I96MwfznK0px4JYql7pSrIB8cn9nNYn4MIm
spoah9ex0gZy4IUd1BRJdr7085ZfRrDeDYKvfhbW+t7QUt+1jr/rMIm60Exx9at6QsyY+IuNvZc8
3yhSu8y9V7nm1VmcQSqEmYOZ4oqT4TOMcNGwxYpMv2Ap4/uHC/zmJ7zXy3oztoN+ClxWj0W5HVeW
2FRhT2SarL3eKZjoBtisrBA+EOz0K6pBLJkqFE0XaMQ9mwijR53MGs3C1ZF/58b0bVC6BaB82WEU
KbXt9m29P9QwunJfQW968YQQOsAA/m+JN2TwzLFbXcpwaa6ZmF+RSNGuiDWLYojUcL7c92gjXX7b
f9PUNp4ZfBumcGkTk2oun0DdLZYmPHpFyBAt0AGgX6MGLFy3r6ewYDYqk/5+MJhjKaIRof6nD6Jz
UOYN+cOfg8w6LuCGlZ0JN3AlBH5b0pE+ILVNnXAoYXXX0Bz9qfVw+LhrV+ATrXPRcwLSMbdeLCsg
IWWdtXcrF8gm4SZUxxhsVtNKqcm43IvM6PU2MVCW+cC1RIRdlWk8OsQoYuMNE4VKwA+tm1jqqC/b
I49AgB7t19P/lpW1E98U2H4cv6L+GOiXpRi+QvnoHd9+eMM7xl0T++4pVkBLNgybRyT9Upo+T//O
J5CDujZKplbFKWuI5ym2ktSoTjRxpD1+Yc6cGgO57kwSqSWyP8VJD91CD/h/8BMOk5avWEnFV7wX
mF51bDz/zmhioCWCUVv85apWzEF+apPYfMETre9LeDE0o04msr9RtoL1o2/6uAtjGmjf1hZR/1F4
sR09aMU6hgQyab9H6qaOuPImKfUwlF492Io21+AZAACeMEKxLpbtUuTXORWBnpaxbo5S3E3V+pcS
kL/rPccok9kOM6vwIt9bXKIUGchQNsbLXZlrfspCUO7k+MK/QChKTGRg9/bHRa8XDk8bHn3zIR2L
q7kyqp1hPihH+7MN3zXGCgzVLryZiwfqG8OlZvlqjHunMg6ktKRENN3ipZf/XFPqmmXeP7aMEdYK
XfQIfvcm65kAy24HYKaMCGJ5RBmn4BjoCQoQrk+YgoG6kvr9EMInlM2xVeCPy3LfH6KUxvRWgS7C
iL2DhbaAJdJ9bEv7s1Tcf3zFOenFX9kpAho3Cp7VI82iXIG8/Jow74BaGD+Xm8sDnefvROKeNBcY
bu/ovutHgoCxwXlz+EiVsbTqUcC29S3HJ/4UesBDzgegOepT1bsI5T065z5TkCRTUyLZ423mD/La
SzIuR4u37LNAT07DPr7yi+V19lrlFdiO88+tQi/b8ayG7Vai8QGla3R+eFjlpIbzhuuIrxJUg3t0
UgSdPe7RbuomWjODO8hItEU1shL3eDiPdGOpptPNMhd1pWbFwXRDphtc5vTV5q6Q7+usb63RTD5F
hxvSsJA7DXL1ZcuilxwVCKSdhJAEnpWbgAN46XIENfHcxPE3SBj8r39L5P3Er0nQEM+B5YZRu2iV
GhDreZ/UjdB0bwztTonZRq3UHDvt0rFRWYF/gSpklCYiJZIvGfdcllTj9uK9f624n1j3Wb8KdPXn
bxtfqXie+tk8WvWVp5z5FJjOsHy+fY0DZkJpLIFnNGUweJSIP2tfnbec32zK+iRceUq6YUUNkoRq
Y1fCQi7wcnjNSaAXZbUDDSQ+lDQrkUnS7vt8jLs3WqLjELoQJOM1SwgNgS9O1jP+f3XnXJABDmjC
Rl66R317wMmyKlUacMkDYXZXEkfY3kwnvuU55kNxH0Aq+6HK0LJtBZB8czSmLDq+FIMEM2he+R2P
o9NG661+cyikh5MmSpHvqnyDxROcypML3tvpgM+JlrkAkNRN2rsf2nRwBbkEAjTMSe3vP7THu2hR
WQkheGQpt7VY2AImCdA3d2395cFhqVZvtHKiwDzwuI1mQYcLPzac2NAROAoONH+RRsB8D5do7Ohz
dg6nPXkHPOShUaHhv0JOYI1iBwjEeejKClHQvf2yNJaub8Zbzi1Gez4giN578TJApPA7bG2hoYBi
cgImjeXoiobjPeqssAUkohn6Vf6ckjccXgGdFmtR6xwPaR1KEU7ubyylRGIvZTCyImYYvo86PtJy
UnuvgocPUp1e9x6mSQT+aai2R9Djkl1MCAaJDzPtIyO+KohOZmL2Fzh5QeGCi5vsgJPuUaQVQM3y
4QdoD9Fx29l3yC9es0oxJTX69urDyQOg9v+daMdEpjslaSyJacHVZfMmYkLqwVDiKIOweuSRLKM5
4cSYZBE9/RUm+SSTEnQkYsEJ7Q3ivbJCbr06sp/Jp7h+UHbi69TJAg+L4WG8v2SwTGjoRmftCN0y
xDJY2f+9sdMNos3KXQNAoT0uZq6FuMIu0thUCcyiyc68aKp/garvQCRqgpCuHOFenf9KITuA+xM3
te0YzP7oFRftXOFOTaRtbyJgqCr0dxa+5t+PlQXsQBmG6Blvx90Fy8mQqwA2XFkly7V8/RTi2Xqr
WeaQ4VlQnsC7xWRSKw7Kjp3kA9OZbHCWAYS34SYo5c2K4nQV181PcgIyMipJQmtjwjnJmxgsGeIz
BAkaV9C/Drkxp0i1nfW7ais8nYv79u9C+HQGtr4RLboWcWVoj4wBZgnb2JrTNXi0C05bsgXoRWae
tIRru7UeEJBMGLKwgWQjdku4XSdMwPZuDom9gj0yE99NTPSZIiUPzUy1hJE1XWUho6K0kXueNzZr
The4GWZ5X26hQTszJbmiKUvNeDV8pzizTIwFzlwx7J1i+UMyaF6Bdqk8s7AMQ+LSoXOlCsLFKnt+
CqyjqDpBFvqhNjzXkhsz7IfIGrXsyfz55jVG3fswzXH/VSMUVmeK0M2Hj1VLlCMCWA1VXJyCG3Dq
Y9OMOqSA1l/QhG5Uy0nf5ZHb8aJevr7oWIKvBuB7CH9KYRtUyi6ISfJIq68FqfkI7A81Ags1omRT
W4+9rYbwBF1mJ4jna8gzghcL4fcDLIg0H307WpBPVejuiYLrFcUij/KGec+l6PXRGhvchPeCnhfm
37gN1k3k7O7e4URPHXM/wR/hwBvESsoTRgi6hiLTN0QZmIqRxoRPQqOHuT7no4907kTvd3MS2WZG
VuKnARp/w1eeCs4ov6gy0KTi0/slmaeuL6DqkJMUf4QX9PVUJ5yakJbju15ZOpSStRRlIz6qP4j9
XWaivqQ2COu6V6bi4Zq++97QOIg/3imx/dJbNXbAwdYyX+cBS5wsRi6zE6VOfzwgu3rXaorOh5YV
kbF/nDXF6LPSt7PkTE3C/bZhDJtdfaFV3tjlOf6pMnFvt6VT+SPnnrN5qhcMypXuTEvC0tw6SSw8
tBASSDXbcC54V6M+qQI7L0nV/JJj/wHejrtF5oJjYswHSnBfw7gmhnQokoE8gOc8I1IvEc5G8+6Q
a6/i5lUDFyllUEXZ2RUMCMIxVOTM6OmbvofIfwLNMGlfZPZC1c3iHDHG/GN35UK31yplyBYtIpPH
Sq3gTrTAv8e0QHTsFOVfj/3HtAIwOgg1DiNbITcZ1FUCZMwNbpJYtfJA/Gq6PKQerPPT28Cc5imN
ChbaqtHHn2U5JA4/r/s7MjhDK0GlJFS8A8pWgjUsrTqNb8PbzRuA6XP4B357co7xOR35I8MIPruB
z4c4nPqx1QcMp8jiXPMyHKKURRaXoWQ729adEVsQTSmSCKGebTVLkpKvIjR/4d8fgl5qEnLjb4xZ
qXbMv0K06NO/Ax5BtJVh0ba0/J+LCybKeMdGM7pRgenQuc6DixbK8k0GZC9/u/kmEafEqlV8Kmuu
49++xuCmJ8409s4KnTfNhS57ZmE86ou/LLRYTx0ZaX9YJNDnSatWHtv1bNxT8vay0QxwC9fWC9Wi
6evh3vpltdRgJ7EUKTCbPufLX9M3qMjUJBjG+manLAcxSMKIlJoYBv2esP1SmiDDWfON1UPBZ+RJ
CTtEaED0UTu7V3ChUsSIQjcHVC/CmnLkSCl/smSc/7DJsuyZo6zpRYEqasM6F6M8FxP/Rr1mxHdu
vvRDyQRgHLCGr1CVl62PWasre6MvUJ2hhqhao+4DDMk28qDB6xTksATfbcgyH7uETu92rIFlf+v4
u/+X2/2tEbmkIy7PnlD0pN4WA81OHlw9GdsXOl3U6hjSfPq86+pu7hzPnwh5u4t9U//K2wTocJ72
AVorDEfcWjwqYohtIX7gDgOPFTtQZ4tWKwr1e4cHInAwgPwTn6fXkByIOjKwyui8PKSU3idmk9tr
vqQrFowvgiHXGKh+yjRr/OzLr/EKwNOSSNPdAba83devTAK2fcZsw5AlP9mS21oGmV3b7lhD1g1a
iI7omkkPeIBLhUrEsypeQeHii6uXjY2Fu2DXKR0si7qr1ExHK1oL0MObmnXnWi9QNfdrjwyUOR8J
n4z5eQFKTPGHi/YTprF7lutmyLTKgtcP0he+CwR3bzT7HG9HRGz8YP+u/d1qAxgGsq2xPqVRt9gE
1Pd60xhQqthbpCsLzHbmecsHk4GNQBR6681OGMGXPtc9ayIx7oerVi7oL6x1ezykpergqLtTIi97
CfzTFL1X65X1HB/4TOHDGnzp3amDZCsV3nzqh2MoiYuop61kkrA6/arhrgabnJn+xgjJYT3RXCZy
CzsDGq4QY58yRSLUAHUszcv60LFc6Imn8pHFsFEP2af3+VTxr2PbugJ5OI8ss1PYQxq/eS+QslNI
Asj3KAbxgR3h4SQU9yE78KqBVllbIrs6ea35SWznswjZ23DQqnUUI+yN01Q5YnSQHpz/DNbpcq8h
yxOjrHyfh6WQpz0kYvXpYKtuI6ZbjPeHW91WITi1uIfBFIJF8G8t9FrJv6g0qIcjYBH4GsN1aCIa
PrUZ6jHSMPQ+6/0Cs0XY9VWVawo8uMM3xwlqi7J3oLNKG4EbalJx7rPoO3V/8tCgBNBkpH8IVZz7
p+uCzVyCVAPduOl1FV1dEi+uBBP1Rpo5d+wBOg7tB5/lFOUebmTTHWYTLgpdu8ltl19Ts0vwFuyP
wg5qVHJ33qD8I/YrtFvFLFQPDg504zrd9xCn7FzwA6/iTKf7tOy4QU2vIK1gEzZeENo7UlEXsUNL
PAo3m2uIp3K6GwuRCJnQrdTYTRicGkZS/CM2ow6s5KZ0G4U308WbfT/Dyf2KODh5kZPgd5SaDFBG
NpIjhl+DjYMGhfgp2JBGpPqQ3uAikqGF1MztGG0uSSxLqwx8/Pqck/lhvdzaUnuIXL5xrOBR75M+
pa85vEenFmXTzM3hw2sb2eO0G+gYY7WZOCvPK6D+3RUKuFM/xPIISQT0V0LvfuzINOJD41KIw/qL
V7A7zv+JrsOEs67nKwggic05wc82+uwdH4PBQJRNm9/lUFPuTGZ8LKDT4TKg4644oRrnulJ7gC4A
WRCwgl70dTmtJ1KtzOBqzlhee/Lw1k78Ia8dl+qrBtc4hxI7Ke5uB2ElW1bf1H7q2JfaTy1gyJru
4iXRenCoySA0JoGfbW7jlgVE8j32IWuLBBMoT0EBIEZxSTTMSLx09pU+uQ7N/bYqxSfVYgSNAp23
a7pyZjMg4iwOAbyHUKuRFKESRCYAboLtH26oU8fE8WU1cb3hS/EJ0rTkMzM5HO4kZsU+aSZvQpzX
VGYA8UqhHybyc8njRAofNMPuAQ8iLDxQUMvxNevkrzv5RO9u0e31xAKOGBXLSF0OC+ApJkdDrOBK
1HAZ68MkAnqlNnwFVBtRSct47TjAmUmU6mPgKCBbAftsy0lbPNOIdXgVa0Cy4hW/2zQqk0DiqH3f
YlMp73gK/JjzNwG+IbF7mdx+3mKAqPTGk8YnvhAKpx7Rq/DQoPENe3MNg6r2Ej3+Bd3Bm1Teh36h
YHCDszpFKLNHyJKHGxFBPbP4IsjDvFcSjggM1PqZhos57Jp0JE9GBaJ6NicSiN41hLaBJla2QraW
PAebKji1RgRFsRRwTXtleAAUbqO2o4kK0ck40V2imIsORaj1sVhtOXEDvKrov4HEwluzi/P0g3WM
/TD+SnJd01MJZ1ZsC65x5WVJoq4Gx9ddEpVuQ/K8CpccLjJzM64Kh6hyA5aTlQ75NuzPjz7McTwG
29H+a0s/Rc004O2qOgpgA42SfT908XcNCHLdzDDm1TkU3gMCIiP+AtaGhmhKjVwwJwAOpwvfEuVa
IKWe1gLQqDSctjgkYrb0ZuAF3rKIHec+rsJAB1aT/QufNLLCxT0LeiMYkKpYmH1f88Z7vOQSjYSG
z00qPFYS+74E59EzUtdF2ZieeecKwuDR3bjN9VedKf6KKrM0XoJ2RtQ5D2NqoG0/PhnETazlJarw
siK+vaedEPryPeiqjUkU7MNSievQT1tEUmmK1D707yT0LPQVq1OqujWOoiXiXox0a8u22yP9ksOf
Aer4hGDQKlxpleZuFDVLsaaRs6D/BN6wRwpXE9refKtUx2/YeNL89upswWv6mXjkyMtgy/oC7uun
ve1FigR6ioG66KIqHk14nSLfhgWiS2mTckyXbR0JUwX6eR5AEMnY6MVDAdQC+dXGfxaIIgQG116F
4TQsVaFM1xOtqz6Q6g/faL57xx0dibUyGnhTcg+KfzNYy4ef2m4HB+4v11FDfTbQqTt44q9aIoyo
uYxNZzJtG0lyyzXyL0eoqaoqNEBid/Cxk30HkkVdOQAOx+2+Sq3OeEF96VSItDvDwhI9qSGFZk2s
SuJJlNNzeOHwZMSJpt96alX93GS4IxODBnXk377dEn2kUHjdwFUyCRUt23fcylCvoPyCWeQ7s9mG
3NqD/U5HVcbGwkZEGedZhYqZkK7nR3Xd7xWPUcufluuC8N3hPXz+KleJyqVtA5xFwx7VAyNVM027
sdy3G1yER6Yoccj1zJbhAogatiL0Dlc2fPJ7ed2qTBQ+/3u4JRL4cHgIUak6PnGRHyjiyyX3wyTq
VKb9FW2TWseivQBA8yAYCRV4CqejO6SNuWjZ33tgaoZyMEeGAt4ay5RcvfQqVRHrL/V0SSglw3fU
lTdgc0EABBduvbEK6dA5yB4XuSmDnNeKvaBhkmTEC1slfUyGauP+gIVoMGG+Bc7T1IdZWAlwZEr5
mJ2IxNcsLQ216RDsZD1ej1iH8tnxbVPIoUpG4xLMZLnX/nKr7cqVvCPx0GilFqtsnbxyOtxLOT6g
kGDf+6Mtivbb3gEOolUnaFzeJRwmg4MCoKeO+JSmQBuUiLozC9ZpnDC+jDcBrDc1N1kIYCeqtRGH
cHkCdFHZoUACmCZWdcW+paqgfjP/SCgxD48Ub9QbqYY9YhU//sQ2gUVXRP86XcAXM+uPyXKVYiCP
KwbNoByc52lDqxhvfb82CWi+xuxKZcp6VX4oERVUU6GQG4qw+GilNMHuDF+jPE+2b+xC4Qulrwh2
IHN/7YRWEvvLCiz8ZVQr7gCQee2RDtZIFB9wubXNooKnrUMnlrpx1aDfjWQwyD6vFq5X6BqLXYsN
MvANtP7QdC0iMr30uq0ZxI4EUQLh7f8J/y7tR2VMD7KWcGv1ck9W1Ru3BfOrEQAN6ZhEGXGSZMsb
flHzS+/QlFoGONS17LUCjQ9GhcLmJKuVcINO0QSgB/HvTa+TkbNaiqsWOHe8Bt54tZ2RVF7s7Wf9
pOV6xKePIuioLMWc+Fss1oWy5GplZ4O+EkBYGlw893Ha2WGhbjEjR8S1ekJ0K4wSIMfX0fwyRUi1
68yuOK7o2u3a427gmdsMJT+puTs8Ohwh1wnCAetipvvpMasChjzfeEYPVM9fSwq9FUUXHQRkHo5B
V2tFuz+Ussj1tRIBDtmEefSSpXOSXXBYR6SfkQBETHlmzTVY8LiMhBYWt9l8Jh612wYETlr8luRu
8xb7zCKvhBU06jvXShue6TuPhTGmdeEheip9Q4xvXLJNLifZ8DYeMUrHt/sCFnfF8pwXbI50MfB3
nnjipIqA3KjQXmMALwmTCH5LOicMkaSKYNaHWwG0ILA7qCS8uGr3fv1B6lhZNweW3UF4MnxD5euY
DT5lTvyAn0FPMO2jqRzMDuCSzzfx9Ss1sWoyZcJ5qZ1oDsn5G/AwmwrIU/G7vOp2mkMDakpooXga
SA7jJ80XeD2kh+dQPQOxU4sMK5UbXkL5wg6fcqNhS8qg7ArmhD+5EEXtMSxaI1KsONyrmpmNWRgx
JArLMzc7mZOezeIdnmg3kThUNNC8VqVp3KMye9Tygivb/SdpWe4X56kvrENjD2sumeCW1GLUVSnf
DZd2uPFoQBCBrD6uXUieuTCNruyMs/w8LQMY+nPZSV7y5OscPbcAEh+RuWbn6mF2SCE2IGNDzIgG
O5oKPrMaubF5d9drT1mjEGNWfX4jAi71USffumv3sJpZ4exndWeSemdjjozsTqTE0aNRE751M+YA
3BWbRIg2MCrGN5Hz80E48AG7tGHuQTF30ik+gt60NnyoXIrUUoZwKRXim0GPGlRAkbYDe4n0RsXg
2o5QBszwxWN1mwRtOttjbO2HekjHz9+BmcdNr3fA+vqD6E4IcO/rgPceF1t+vTaxQMIH+FvGzhDq
icb77jZdAR00PdbnTI/d2GbKQFYcvG0q6ZdNrLvV1C9PpfqCTfUahuwrj2MDSLyJiiERXMP4SoP7
WfqT2M0UjVQBR/5Ly7AcuE+iJRx1kv90/ADP6SBo3V+G5em7b50Rww9oDamqYNZ3WViAfIAijUfH
y8hqF3N1CkHSm/OdH8Mh7ncMOp/PJQ0VkJGquXulwdy9RnQyJgBBnTisqgE0nYqn9FumFHjGgNcx
D471UFSnCtQ16u1s0z/xQ8Leiw8JTk/fE8RGADf5wO+9mcp0vPQ1MLw4uwT85N7GoAEO347ZTd9t
QL8fEz+MLosb3N1FqiiAbHGVGrINq+g7ZvXVugCfuqxWmuIbExoR9AJPMW1KdJFbtcGbKPsy04Y6
ccuecfE/hLmtfcxw0Kxo5tHINJEDWnkAm7+OoV8agpixp2+EhaWeO6cmFnWzYo6KnNs+8MH2Q1EV
gTuFxY68jekM4gK2UQzkVdBXYTZKGV8jPAPbbt0VIsPoPK1DoQfDPsL+hEmlbxRIoNDZGdTW+CUM
1UGmr8JN3QS7IDiHekkzFxbiaXEXA+5AfpdYiWBzrQ/x3jsbIRsLWwdjJFHh0cmdDX7NpWAgoo60
AjUkoWtjrAYeDZju1OZpMttS8G/m9hWWUzR+oJsXKCPeb/SyeTMfj9Vk1fSVZKSllI6V1ChnLWdN
VgE9csprhGp9tTqws1A5i/YCwemyEgzBkWhWxS7hN98ZFC8PosTQEqQ33FY6/H7UA4kQLeHK02ZL
kuAinUzcqXdfHImeu3x5zhlWy4wKJrdpRNu4X7vF7PguH9pr77vIq/l1h3i384XbBXCnJDpPD69K
1EC+hWfSdwpobLDYpV8QJJUOzAx9uY6S6REFqCN+IjvWPsDbRjUjlsDerYg+V9TsvjJxpYks8F+9
7ka1q4IJfO2EJmxPrIozmCQi7p3PMdnbBexQFD7/OCw7siSusxqgnWmXVa23hDxNfoJ6Qs2i0OI5
U2eWa9fCOjgHPuOYwnnYLEXygU+zgAYpx/qG7lzGVFguaOHi11YwuScw4NYaV0ThJtc8JpmauZzj
qBqRkB58pvXNm4zA+LHqATOyBtjtPd2wXNjyOR4eX9ccgdWyNgkkA54MpO2/uAtM7Gk5x43ekrlL
AG+30QCx/4en+iFfv5G8wsnO8xOHxDAapgae4DjvWJk5M0rWKFYCJDPuZGMrDfHWta5/fPjrdnNF
S0wMteXiGTnfCm0YPGoXks4zFcwsfIBWkqvYadv6VP6akaGnyRblLs/b5YfG8tJlZkiptxpxUsFQ
0tSyZ/a0zKZg0xkeT2+t6ykW75OIsMeFteQ6S9T4eI/+g6QgXSLvn8w93sBCKdMFYobVhiMpyQTn
9Aqd56mEv1sK3eZFae5+PSlm/hCvUnAWuFeg8Y/Ir8yby4HclTJL7bYXLlLDM4pqSUIqgHabqIwB
5Slr3Mi8yn9KpRrWkZ3XQmvy1xaCD0b4Q82RA29c/GtG8Q9ZYN5z9Ui71SVG/2irTTjldhNEpGD5
Dbk2ilXwhWy5CUaxNm4FmGTEJCSXjOn3nCTMCvGCb9Qzc6gnpCCHwN78PvPe/SBdeTFxPcF7Cnpn
oPOXF9bRWRpPQETEOTT+piN5pQCKNrzu8x/9r2MPv/Jp8Z7zKpzaRxyfluv9Myk/u+b42wf3nEAG
wL4kjmCrfTqA8Ef8/2MA6ux41GpyVtviIYbaJpedkr/WCDMYL7DVpabqW6omwTNvAGbYEVOJ2MU+
vdk6D0v2xQZk+cMec9fMa9bItpAIuFl3qudttCnVbgb+EMwTzyeSrNCJ+G1asSs4B9BuUFwAdonT
kdYO+neoUG6eih/h6Dp0VOqhEnv7krrLLPjgX+o+OrpePcZRJMXe5RfrdjCoVCwam3Dv20r+lNK0
T0ldjEt49oC/VUXW6BP2a7X9+B0GL2Wk93JqG+C29yWM20wnJ9dn/Mt2ouCXmZ6InUu/RzWnaZci
YN+30dpXEdNpaE9lUqoil/Kd379N2dwhfa7vRbh4SOb6tx+uVbkUhiP8BY8TEYvO20NWerO/HXKr
FwFQz63z9+czuvmhTZ5jAHNwvzX1Z9O+OYkaEqrtDZLUL2oMR+Laki3BUV7Z1j8L3pausOzlQPCO
eNE6umgXSFnd4ezHk6cBTVBS1aJsgQRiF4PUicIGP+fQz3nT4NeVvbaO/LCm0mxq0pgqNMGGqATx
8S3HwzgW0KUlHqtoRQZbEuyQYXY2HlULwpfQTkKSiHu55HmM8PpMoagnV0bTamNf2WAOj1X2mJkH
f1MoH5Q0bn9o5SQYyaDFIsdit1GU9OSqFPAo3H+xx5I/vEFyVW9sQIZvDGsDhzlu75my6XWmch3j
0PjLzuEp1tV5BPsdEHESdGuBIzjA8f49u39ZWx5IK4UC52gMVhwhRUu/YhpCr7DMGTh9k6kii6Du
xPxbayeVpfH8+u1dKavymwpEnkhbW5JeyqhFmn55oJbltGjcHGJKVUCtASXB2DAWBKs+sIPNDLmQ
LJavJA+Hs1mnF3wr+DoIawl9XIX13VAo4dJgCIVmOHgKQWJKRYPUCyewgzsmfF3333P8JaRBXuPr
Qciv/ithZAXDoCtkivFuYWBvGaBqfsF/hwp6dMq0OoSrDUcGEkRpzMeCzX8Ay7zmqH5iLKYgj6lM
x1/Di+kUwVjZNrn2Fo7wEzqWJznjmKavFoLLzItWAWwoGjOpQN2T2xouQ8QMbqon2mb7I+AVNmGB
zSCDBsmvJsPaKs8Ac5Yk1w3ZhMDqLHIcNu/AWuzyy7/eZ28UnFGR/4JMhAsA1yARXDPw9a8VPtKA
YMGXxZ4tCljctYvztmH4qnSIgaWg2KrJlUz3FVPRDLTgIKoGeu5KKFCNSg7aQuswIreQbodYc4QS
hXeu60j7svna2DQ2iVpjtilry/QbNEL3QEIY9KOYnA6dsGDrHOu7BkCO4Ay7GQCILUPQoICjO11x
x6iPvw75RC80XxEDDPJRMPGCezoiGe8IWAImZWICxnsJGleEvyZvs9m1VcHmm+C4IFOxGXLDyHN8
v1QFsQGFMOKuhU6cYUJtyuT7JL6JTYwbIEcfPrP9fBRbPaEpZ1HLS4ql4tEf3oHLIeTcUVyHmgyK
/o2ozWJCtAQ816RheAJHJ+PH3BVUGFVFXzYR93kjwP8Dy5KNSDNEzWv0wexeF1i2uuy2Lrd7uJRK
1Jb4ulwuPZqp5RdEEuBzrML0JGu+xSb82476cab5UQCaOIA2zKShogHfLiAWyfLRfoXWf5O80vsh
dvA6LR5tDSKJ+CO9FgdMhuRX8pgRFqyjzNyYIJaDZVpFXgvjBD07hsYQMu9IMoZh0LB9AOrMIFek
NIwN+HlcnOJKiOJzc2cPBUQoyACOLxC8K970fpnVartY49vN1QpIx0eH7b7yXg1oFiAvJIXNOF3o
SyQ1BEu5hip+ZouFGGXjidL8OdxRI9Xl5+qI1r3k8x3SyamloxLwsGk+0IXBj+IvRIXhRIR2RJ7E
LrL5AsyF4a2LVC2XgwUGVO4Mfy6ivPNWynleqnOeKMgjr+kC7oU9IxLVecyrDQ0csIWTtoPBCijl
DWtW8PSapVjTi9gYl6mtpl5nnKTngx99cmNCNV4YmNzdvd5nsxqt1XYVBGHm20T51jG7PshvOHjQ
JPfhScKbPAaVAdJ1/upOnPIVmYlDki8iUjj60LW81rFYbNl9YCtmVkiUXsiOUVsFb5z5m3dGlTuW
mp+1YUPcJwyYo0FCiKAX6liSnpNd+u6s6E82rcgQ5AY1NA8w0GBfyXOp0w2/rfWl32T7zNOoSSxx
bjdQbI0Ap/tb3KZYtrNQYsiwyd0/6Q66+J8JjpIO9dSukAVwj2PAt6UM9Ixeirltp3FbmtuGciJl
cTlVidwqOVu/lX2i7YA6YsbYCN3NE6l86pAUfLa4W53ITp4tnajlHWFhe4AVPI6D9YnURi9fthyI
kyh72o8O8GqZuc3K/KZYXobBs17NiyON2qfcgHBryg4MvGRmPsKsT5F/g8ztjJWHYT/Nw07u9QnH
OdxgFx5grGsxV+SbhzoTQJDo3nuDwMR4fC1PQYkm1Me3PV8L4qn16qRDAH7Mdyu63oM010WurXpE
aW9a9SqQow2Pk0LDIEfXjke0rJJZxIbena6YhS4OZH09a73ot8+dhxuApcuZ8+VMEKLvrcfg/z8V
tWwP7n0ukWb0s37ZeOIdEcGXXHE6TGKQ2iFIu453KgtEKWAEVyySswpuEEI/J9BpN94R+In3rjuU
efaEcBKqO0qV+KEXLd3fkXcI0gg8BjLrZHBmWnoMeZAjeaB3iNiB7QG2B1IAXtyFR7SNDxDOPiPz
fvx61XPdT2vhUAPfuRYenS8INLQ+cbf25AizYdWVcKuWdkCvFD5BCJcN3nT9UcasQFVxTkS8kHmd
95x3PNB4LkMreIE27P+ExWtHJoEnSXPmk9EKx4+4E0IngeIAGUF0PYEIMX+Zwpy16R9ALEaZwMEy
OCYA40vBX/GxXYx3b++290SiZgrL0PK+RP5+H9X3L3cQcY/yyFcKh9t1fgU+IM0k0GSXupytF2Dz
DV8jW4EzGg2SmztJCpyKSx746Pi+3xS5GcJxgy1f20yLjpGZFnT2SoAZbp6s0k1Fj/Z83HQoUujH
//pdngKHeG/tvyaDy2/ebi4mzI80kOQuOmTGQHywwXsPbfe6FbkNVVdYwuV6j801ovgQHBkshMKe
PQJ9XYEPR8Lz6UOubC2m1U+AZ+GV6NJnkCb3kZRV+Qh10G2QdATK/TeawtsI/S3aBgu0xOuEQPlZ
AuGVRr9wnu8NKH7e+tGmj99T5pU34u9xlw/4m/qB/WuSqUAhCmjmDQ+XOIU6YU6KvOhj2gl4nXgi
pEE9JaBqGGtyTXT47gSkUIyLHJmlskQ9YVYX4Qk604ErXe6SS93xtmX86EzSNLE1skzXnLVdyOx0
gSxVcLsKClUKWXOrFDGEtM3qTvmEgRCNcT3APzj+5GOyYJwO5/Tl2000LPQIteDt9Q2bnl55JaeL
wNjYHEjryqXFDI9Avl7fuYmne0vVE7cRcbqHJHnfntQkCdBzKTo4RQ7pazyoV23L7JNJRAgZOXMX
G1gh/JoWAvu8a8xhqdzWepYcQohZMz4QMBzHWAdOu86udEuG/W6sgcVX88Dy/jemdagD9mFAcn+5
0mjt6ybMMeSF8ceQ7RtA3e1UdXbkq41UJGLumpp/qWtccw6L9FeJsxc16PEGeHiQ6+qavoF8jRt9
58xflHOhf/2xpf3tcPhMmsp3RzhetkKyhmFDsRtIFRUDT5X70OibF7vxoOfaPIRB6FOciHd/UF6z
jONtQkJkNl1DnpwjXmN7bWrOZWUJpqMpbabbKPx3k/Ph1S6IrpNQuTZANUyzqI3fLnzTfqvOhbGu
USdOlb9YtrxQf8ygcuy4EmLMkgb+tyt9ovVrPi4rOLc9Zbsmbqwf/NfFyn4HaNm4PMr/Bo9LCgdg
giBdghNJJLQY4vnKWnWDCG+PUKFTJekCRxo/bLUYebqCLlWLsBHdv/ErACTBdw9hHOG3bfNor+Oz
/a5BDmr/iSwk8CDDYyGk01BichGibMeCQIDDyiDpYfGljhJA3D8xNbHq1UJ+6lzFLXme+pF1XEEG
S7CESERT9MzHKvBOXgIquI6tdGDnoUdTWCFCY5J7vt4GJWTERdekWhYoiDbX82hcthJekrU6KOS7
i1U++G7G6qEIvA5/H9ESRRoyvgmd7cRzrOSAaqCb6TJ+1+Jm/ulPh/rwrF+T9DETZz/UdRSLnjgE
WnphzACBj9OHwP4JWmps7OqTM5A4dfoOpH26MXrxdGICxNbqZmfqxW/e1Nh7gq2IYE9aD1VUAUZW
yEYnemhz0H5vkoMYKqLju58AUIf/Ee09hNmHLZ24HOdOLYtV588M6y/WSCQtm3p8UYG7pdngTyU5
mREX8N8ytdMn0iIE0R1IQb6d4Gzs3rvGFksBydUfs0BjzlzqTcKChl6WrkqTinF73irZtbZNoT1j
84qSBYZqP0XI06o0FpQ+NM3MPzicSe13WrW3evChLdd10WeHcp94xImv8IfUgfUEeCDKCQTOmx4f
xjpoBxY5XVlEg+FpAcICqxslj5PfuBtjgem9V04DYwLObjxS5oRzb5t0Walj1mtVOEEkb/zcAwBF
x2k+I2rSdHGUxRPiVY/X7BwhEJB9NsFamMCB5oa3kVdWevEz/KxZAajjDKpXsqDpzpSAbC+TDQ36
Da7zRULUBvVtFrO5J5SfyQZHDLMESeJ+CQwgsAMvjVRqEmB1vuyfItRa5rzwvGrYWDOw74oapGmS
wAVk6+iOFwmTFl69POJSs4QQ4pm5f6cuuo+gIQeaZOqrA7GZC260MYvFcIMByGFYvYGIndnH582w
6sKkTPeR6JttTJTJyheSTaK67opjB6ryBXzVy5qoguU3qcphbO4lv22Dlue9MkvxMihUpDp81L1x
dBZxgqKAO+X215KbKLm3T7F40YVShZrSCQSobdnlzbAfMr4kkDwdgk8SCSgoJE5V0wleMRTVrnAo
dnPxMRe7JDdFU7jTGDuVgUvtfsN3Ht5C5FlBeOIpJpXWjeV609mB3Vh4oi2yDIoemRpfhik/iVAK
l2bh9yEPgxFZhpykl0WBjMUW8ziK1K8AFe0sOtsAJezWVpRz9uuiCwGWUoQTcFcmweG/l8oF82PO
Lot/W9Ba/Zys+Iky/mjcBPdTPM5de2sUsqglAUrd452i6FnczMtDLKqIJ0IsMcU/0e66/DmJCtnD
WUDgx1zqSw3fkHbWsYUAeWmdCz4rKiKA3fvGSjxwzxe+bTsMsm9RbkT7qWzEs++KmwlUUV+F9ABp
ZMQxvfgwDHET8gNImGOQvJcuPdPm7ffc62daqpSDFRdbqziI0G2SPUWyYw0ZjuzSaOXcdlPJFqty
m0ji8MS0wV1mLEbXwqbW7IBT7fA+vVrGdnOrc8Ntdkt7sob4/vFp3uK1tskuFXlmS636qMlTK0s3
LEPvM0A4XFxVtVuWbeWCOxKjCRDpdXz0QEMT4jvU82YOjAi2ifgLVEPW/xCvdbF/nwiI2wfyZDTQ
Jg8uVs7qt79ON1JkSPucZHexR5TQZrzA9O9dvcTCmf3s3yJX5sbe7tMKmpnPoWNS9jDMTbHQnV52
Ng1Bwri2bDg8O/akpvy+S3LeQ72XSzCCeouPmTcLztv3/sCQV9E2T9MBEqtvJT7OiFohiHgXSldA
0pqGe6muYk09as+1wFqKSoyVaFXC/gOAsT2G7LAg8l91qAfzHqFoZgz09I+b+jTfiAB+u436h/ea
KWnJT45OjNMgAg8+Z9qj0Zxeo6FJQC72dXGnEnILSvMGd1213SqkWdeunQDNsdyI2IVoRgB4Ad+/
qFudwWopXm5DMGir58/TUOuISK6+93Ezz0xfDD1VoK2HCTXI2twqL/OThVyYDdYovUahCWqWfJ7N
OxG1STLuRPZWDqLgE5MH9aU7vO6fb8wLQEMg4/8xSPDTneQUW7J96MRHZsxrIKjY9jqemFDxWksd
ulIQGSa244UWE6Q5JCW5gfHTdMnIN91UPhZSvIMa5ueZk3u52hW+zz+rZ9YYgKxmEXDG6qPyNq2v
O/A0y5Kaxo0OgOXs1TCjPsoBBgrVfDcCIsyzqr0ARHax6fU4z3Oz8qi30060qe9wZ3hfP44PzZam
/CHRe6sOWCjkX7dZhGvn5zm1rpVDYz3Fuxgv/8Gqo5NrbDciC9OlTZ3NtZmWWrfH1GtsSUuZURTH
gXrxtFsEO30aeV3krK74ywAasI/QYlCP6sGvelCx1q/s2MAoM0U4C3IBKjVuHeXfB8D79JnWD3t0
6WsxY107X2R7Czb/yN3p5hlXSImtNnbJ1D81HrVrnGI2RD/Q2RqFY4JQx88IPa7FHaSCkcYinZdS
8j4qhTrLMBbBq+widhrwo0qZI0LtQpZ8iz98DPHfvx4sszpB9seRjLLio3k4yegHURye0/0mpqU9
GDV6Ir9DJxECvw7CImJrjfLCE0xZZ8NRuexQ7IrsURl3GK3R5aPLA1tX1zCrFq8lgSrCWOQYy/ne
i0KHQM7BoolH0vhRk2kGl88Q+3IfTRdP9AJVqDZgAOzd0aMM9PkmV87n+f/HJU+3uyFkNBmfr+YG
3XA0HVAats+ugFvaEN79qcPRWvzEuT/dmeWCVzUkXcWCe3vj4EczViOVFiTGdkOgBrQQCc2+Uqav
ebJER6ufKy9GXVQQgsv1Ea6b5lSHp/FXHiQwXRbqzoFiG+f7vvUOfdtKf9YS9/MGsHJdJVW1dmdK
7iJmvcb3nTB6JeVBdIxAivGeVcQv3SHjDHL5nuD0NNCYMDzjnGGIOL66ivfRWSzlJSZOdWIsDqwS
SxVjBL+XngZWa6QYnuU2bVTEqsJ6+FvvVudZm7+15c7jOXxFWm80Lipwcj5WzmEV9++xPRWRgJcA
6xwU56TmIBReykDs/iys2n8MbzC6xUq7XX1mXK4pAN4q0Qrz93xhrcLbAJEU7qHdkNt1ganxAf3W
QAsr56zgkyS0smDGq4Rgj3vGw3WBjf5eYwN0r4A94OapiGLPdaYFxmxJcY66n9FWDtubtuSZ/VRt
45SWN4+ZHwMEek1LkreEElOLZtwLOBPbDOW2jJfBKsKcDXh2WPBUHFzxQfWbSeDVreZY6sPLntpA
wbFHnXvUEZHRJUMek0yleSEdq5uG+q8P3L+s+e9yCVf+nn/zNHaIvWRnIrT1L6dZ67jSGX18d14w
4jwZw0i2h8q/TytZQuNFI1b3of5tWR4AhCWMe8x5876pRJ05JBYdQrsHfvovsuFSvc0GMlaFU3pI
SMCBSmicWVFlfIRZVZx4MkWX0lyn6bTEvLv8zPERMOmR+8GP+P3A9HPlnLzDm8aeoBGtCD5IWyhP
/wEDvGfauzceH3OrCRFDWfIkMSSQ2UhqrLemmTPJ59MqxANkjMRtsuHDkC7Zo6ukqDmQXEfiHlUX
iXAuXuK6jMtnmg58/ep84qInfoTuUPDI5s1HeC00VLeu46oa4DTgPXwICq59zZUJ6CBheClARBTm
pyGRJK+9M6CaF8tx7d6Qeyoto5twE//l5N21aF1pbgL7S6Pe5nnCFKfK6OdHbgjfYDxT5tWr+vhL
ZdEdOU5G3bHhNbMBm6rWog98ZbqofUURhwrUTO9qcxg46sJvmVdR+g9l/9fwKhZRvYfs7rbnMBG6
GwFv6tDtK6NeI8/mjWdEdtoYRkXHQ568cIZlg9NT34zhvdYombtcSTSpCie37A64/86i14K06bGZ
Nvw5C3pV/6wMT82ROT/JyKAZpew+jtRIFsp9jwUPcGolD7cXDxx06qDQwviGzGCyLMVA3G/eTjHy
UzOXcURCN/kkpdmmtcQyPhwCRi2UoWtYNVmdMUI22AY+f0b0y3AGqRQxqtgzBbKfUXBTUN5bYoH+
seby6hKElBiF6W2W9Tx51y1780a1P45GjmB/YKkiDJBeRjmThttf7BRXRX232IMEmGYR69I1chP5
aVFT4MkXlCLAgBUhWa/+IwDzt3SKkY0dOThtZ0miyyhTHTrEyaRMmXYbLq32T41sfrI21EPLTxeK
0GWi/6PYG7Zqe5h2gNK7U2w5vho2+O6Gdc26MAdz6MThfjOJSOcqZc6cBGIrRlVm2yVCA+r0nbaO
klaZR0dHP9topxlRQIeooTvqx5PcHF+J47sr+PeTtrumGKx7Y2h7SvPCOG/idjB3Lq7zh4r86PxP
/CX43ColrAD/ZwONwTJ5RwPms5Yv74lDSTA2zDZ8Dn0QBYUfd+aKAHKwhr2/mtU52VCCN4a3FY1c
L43hctTDvmUci35QnJZVjzJk0HKJfFjtZO8nrhs1j/sxbG3HEckaBDjWHiifMheAoIQJJA6KzDeS
NnWbIKruXndYKyv/P48jfZig9EOHh0gokrE5ewDu0Pb+4F2pOEVduusMi07rRcoNDtiGzhIfcyEw
sSKLDXmPuYouyjgg61YQX/i/EaDtLgFvffWlCtvTrw5RC/tpQ2DFDXYVOLxlY9k7pLE2CnOTMma/
DIK6Bcy0cblSg089w0vD3fz6fzPPUzrOjjD+jTY+lPJZ1vB4UuxZJsDCTw2ksznPri8rkWdaQ5Z/
ntmiX9WVmV29EHRDRVU2z+mXayNcESk7tuFALIKmoW/KKEDMRGy6XiUqfxL6ZtkppGNUCg8vMlp0
mJsXEVguaU/EapGVChzH5hkMIXeZtGRXZLG2swzRr4OIOt87mnmyiZ/zKFGbMHQqQlGMtlf43UR4
ZoRkrcwQ56aPRwnAIZpSvysfr5tjRlySVixBN5saaFwPQsBWgzVnA2sF0B1JsPoOMBurp1JcZVvW
9ps8GESH95iadkK/+oPXy4n6yo+it17+TaNxhbEgNe1BDH3ktI6r2oKTiuCgFJHItkSHbHSwl6+5
4uirzXRYXasFs/NbIEm7Kr5IGYl1TzCwBBU4GYxPIClyDwISmYN+P39/c69fxyelsml+L9CoSbV0
K9jzrAo2n7UXYsi6EhvzsdgK27c9x2bUUjsUJw/ZXQYXktIQGEfyrioq6aAEmADCaQPDfCIz2Iyt
dyWp2SuihkNYJ5qAWi393CFKckbkQOzZ2d1rnl2S0mdibzV/YF3FkSUKWA+XUfKMjo39jgdL79iL
tjSsiEbCXHkQ2/Vg7FT+Z8/Hsqs4/gngfvOBc0wT6tV9E9aE3pYJ0Mfjitl+NepT/OQZZj2TojJl
uv/hgZyoVORH9pWfkwmixO9buxYzjHV2dbEyma3WtebeJ+PX1dkGm9A89KwOfgfyWhDYctP8F3+H
x4ii3LhcsQbj+thzwnuccmCxBdqiHekxL6hl+4qe8/S5uDFCpiaQlBfSYfEeECzuZJJbCje/l/s9
4DpuGro9zBNl6KE1PdlU4cD3A9KD6wwsfTFlg8Pg8GsWNkMQPxtg7L9C34knCc2Jb+BgRrQs06VK
j7l5MO7fPO4ge3CPja6JWfoRagL4voVZ+vMalb03chtN20SGLenG7uS5WvdT9VL/dg3v+1BrkbkU
KoWb8NaLRfx8LL2S7x27ibK0arZbaSPwkri6KwbhdtrHg03Bn+LSmAciTSXlsZkR9+lgMnRLhx2w
TeZClixwv11AS9faNnY8S+j9IY3Ml+Pp4fLqXhIdegMbRyn8WL9d1wMnmJPLDkwVhF6seP8X0Bw7
nJypVcQdUz2tz/iaHBXCtkVkZS5CTZop+hWEyR3z4sijmh5D126azsBDaB+SEqY3lmLvLgwVR39m
uYx7EAEsWTrv4+kZd6QfFk1iywGRd4syANSZnKbmaVCwGhZOUWpUArdW/Be9fEDWWz37uOQMgHij
CIRdQu4uk2huylZNJ/hYvG1P93rk0pxy2oTnpQy+7r9361/WaA0YNeLTjdpCZf7A4groK5cv7nFO
wGb7vj1z6L+U2UzrWIjqpjtGPzqdlex5A62WprjzGW7mKgrZlncMOc5sVGrNF18/KmKArCKkEwAC
mNunlr1hZYDQv+GoDATyLJ8WZ8TVckXvS0sKH0ycmKdg8f1aiVFBDo81cWQ1k5HQpe2MRhLOniy8
P84I2pU++dAYBiISIL9g71sSCyR45KJYDdgysMmrWHMsggnsAciZjICSfjBHjoFvynoO5NaM4Ve1
+73G5VAPc0YJxaOUbl+4IVQhnMuMeRW2UZ/q/IQM4+6rub0SQz9bRVRQXEwqOnlzn1z5oVk0CIkO
ZlK4pM0i0G+wJSfKDUGboUxilEPHARaILbqjvMPRHnnSxU+afKYjlu2BTkn3u6FAxP+aIiI5/dCY
pRuDDEwsZcf+ipgb26r2VipyHtTLaM+nx1QICzzELer2L38nEhwN+yJqK9OKkKXzaEMu2FfQUWhD
b14fRFZmk2xlP11TxV2moxIm0njjUBYxorSh39QvGHEVN4mIce5nfXFRrVyXEe+xTDKmyh9e5nuM
5MYUKaV0caMUcuLp7Jj81jTsi+9zIIuhAhK6MSf0EHXxp8M6b+CmfS0SAqVCP5JchVzm5VCVGRH4
td8P93TQ2Hv0z7PKtF8dJG1u0hI6Za2L7JavxwivFGqvquJjIUF2HccaYMMu5cm+0gikDTTohwnF
y7y3SGLITAesTpcw0OPJ7IUU+0PhEvCk6la3jRhxBFzJLCETegJteX2I8JBMZtIoNU+DqgKrEh8P
4heltQsuAEkJH9UkOFr+dOhyKoVUBW/S94LacAgTjta7j+LSXdJPec91t2LjM/tcJr3OoC1OMLlC
BR8TgUU/TUr6uIhDGgzPNanhtl85hlg/AJosRkfJJ7EgJbR/mUo3pe2j+9FqlvgSi+8pqlX8qNtR
eCko22Fo8RC9GbbczifVKZkOQsnowd1nvEgeGv/F8QOeesgH4pyJI7k3ckSegB1MW0fjOKQB3KFj
U5wSSE9RXj9KgLVshVqEZ+JdFNSfEsrhWVCM9G0L6BvxivoZho3JeFMCW4f3GGvtGoh7aeEhURjH
A7qIjLaRXqhRdYK3tgibxtCnfGUis5PNhgX6NDnsoLz/gwj3dnTtsPDhfNDoZYxIXTt2GB+fntfY
KV4uDqO8eNBj54B1v03MKFcpeFIfR4Z5i4eGiuZjRnrkwSh66s+KiKJi/C0OD6J8kAGQAZuCiT7O
A3qtuzrbhzY1dBYL7+Z5qXoTjuQXTvjxy1cqs3sC3agnEGhzHY07f92juS/EUevHeq7XcHjK2bGh
LbxGebHt3m1bLT7MDiFzLbUPYlTQhWprK74gXTo4+4Fuvs2A9V5ZJDZ5HGIDgamVT6Tj56C8yiqm
GYAFdC49EJKKFevk7ykVACagvyYQWfZeD4HljfNeRJd4HVRR+xecxzDDfno1kfF4MdYuR7wXMlG0
8INeB2aw7l0L7ijbZ8UZngkWu4zLQ+YmTnL/i5sOV1gL1vmvtjXi/UF0khQhFwcEqv/BVCM1DLNZ
OJ+1FksMHORBqJ3bl2h5nGU8wKSVM8eunhi1PRCl/mHcpqpYKzRzpA5678mU98jx6KvOae2rigYX
hP4EoUG6dcJ4b9eaKYT2q5tAel+DINlTQgAUYL7NXZRf1sq/LA0l9UHzt3PaCmaiPf9A6WvB67Or
HtihlaCdciFW8KLoegr3sBJFbrZKvNQRi4NfyMM2A9zp782oEmsnSdpmRZeXbU/ESohLem9+ONEu
kHQ5zPsDLSY12xt731xdgTb320G6AlSIhiu/8wmM7KUIwmEkBrdd66iQtDrExBVMHhfYnZ+AjrTZ
OyuKWfGAFJ+Cmc3aAoG3DTEKD1fckavhluNVP4+5YDLHjAjmFakbDynnenlvo7KLUevpO8dLYpz6
cEKfThcS1JLld9hPPShayYwMS04JxEok379YrjF0WGBKx+3c177poUN5S0LsPejA5Pqx/tuUiPMn
reEHjyFs0UioDXjPcWdq6fzjhQPpdcSrViV6iiHr4se+/qSe0l04Gq9GEJQq0XPvmTqk+BKFo8VR
sZ79/LmIZg2wro5deKR7lvfcLsLniGdu4QqxGYcQhgq4REtcn0/XZOKHsZ6JOfBVn9/dW4/dc/yG
fSvCel8Nd8A51HqXxgeHorjtmNkMBhsU1ryl08vaewxqV2gZblxRMl+J3R08rk7F6OqNF586qRrc
OAnLLjw3uU91OdniCT6TSiDS3BxAU03dXAEb3C8ggDo6rwsvCdxGjia30UA0FsdCcPameB0wsLTU
F6bnszQanquQmTNUmmIVDcZraIJeEUPhyIupiAqr2TJAJbtDZGv2NoyCpxZ6ByX1pqV36hlZn/eG
5RqDGawRYwhFcAvQD/Bzesk6pWvoZTBhRkKX7tNQv+rMQ4iQt/LPXZMAYeFeNkEjw6iHWY+gkpfl
eE/QPVibJSDwpmYSQ+tNVA9w3MEgsFu6PDhGw6PyEtKpjyFmiV8GSt0CNqWLXil/oYriX9fCCDLB
RjnVu5jyDFU36JaqwIogisAx5mEwG9oaAZNJ8IMGGCAoFpl9pDbHtnpHyTTFFwDFHbbUE1EB/GdN
j634mp/awyd1zqRZrwckzVsE45x9dtfJnrt63VSMlKKSy08F3jsvqSscG3AoeQyyk866lGRYAXaR
ow4dr1UA3Pk/1c6b5S5K1CCDiCMwm7dHLBfdPonx9nMINEU2m1Ocl1WyvFZNOI82QtX2YMzc6b8d
OH4///BMyYmwfD/FGqnVP2BLCdSkwBdGsBeIl3rlFYwOAOPd5W8Y2n62Q2SAeyOZoIXcjbtbIlDv
aacBweaUO2xQD1CbRZj/VXiUtkugEzzrWKRanaED4F465Pq0oTPO1Mx4Di1P+kMelJeu2Ys/tuyZ
MOdxXjcmHitYdOyRLYh9+LwwJMKF9O38qR48pvAwVsEKhNQJ6jPlHF8HQp/jPtZ+ZFwODB4njgxc
wegZLW3seH7gFNAg+BsPfNxFJzgcrp6cBW8+cpkUP+uVdJYRl/rbEEG06jcfqpbGE2qeLPQhlvho
Wav/rS7Q8tg7B1GMR1z2OUaZGJv86wCOSPtbBZv9dRcxjgZmPSK4SE88eIleK2pKnmg/FVK2PCzH
QRtbMtto6EZiQdQjgkr1KMQ0JzJ/EPkkHw2d4cs0tYB4xhDuxU0BDsLQrGhLP7uKlJSIZ58K1/3+
Eg9BzJbTvRuhWn7GPv+kRfsC7neqwdlDviwl6vnzNWMEwAjcKtl6ueDVXY49qO45sMOx/WqqF9AB
62GB9ekhRNygWeMO5Fe65eomBT5Hs6gB/D3ft0Y378/xtdFKms6gevVtGuhkYymNISvKJi0QCt1n
5c6KCg+EPze4XEgempHXCHWSdcZcyGL1MGLP2eNu+E1KbOEmGxNSQpcq1LZFdGJgbygnqBdDDjcg
6CtELymnacvbW8YDQ9I3w6B96nCd5Nb/9aDwurMFCajyzaWKs10NpAoqkRa0xLD78fHR10aLiYLV
f/hFo+LZXjbMOEuFdIccQYYcUg3uYpbD2CcJQGHzaCUShhct9kNwvwLfx9R8GXnnMKVczoipnd0Z
gIEdd/g6GgjbGQyeoO0K81rfGq3qxrNaLfS7pLYNxEiOXS6TWy/TQd6qWYZwVLD8CmeEe5ZBB3iE
FWwiEPwcvbc2qNYj/pJFlyYfcEAVi+meuilbOHTJJZR5b0xm7ts+5+IFTdf+SsAoWS1YSYaCKrk4
zBnRo5CKk439epVVM8HXTOXJe13VAz+cQXJsjDgeMG5gTf6pNcETnWUaLWeH1eT4lcal3o28XqcX
aw4lB8y/Nz+FAXEOmmJzUdaYn9M/wxcz11H34WErqUn32XERSe1/akTu5/GJKOUTwSyw1KoO+Hx8
RrLoUQyukRrJMnuXmicH8tiLt/hSnMg4IaqG2IV1NLXL8jSlH2bz+aOATiWk7YiMrHS85QnBwF9v
A0+IfMdZZkesRbYLCTi7ubQpq4d6f7ptvAMcupBKS0WaFiTIiheyjAVw00BERHMj+1JewSpIidHf
Fuk4yei998PAqa+lH6Q28OXt7+hd24pCZMO+YHDRRW9ZaDcBJlpPEbMc6gPZjEiFuosgHlfn7//S
7hG/vCJOkbIyt0hBzp3uENqLujCBqVi1TNlFIaArNFCHLdar5ES8AbFIwduqIxME9s6wNrC9G3p4
TJszru1YJVkhwYQvhSY41OkUkKx8XHRtMmcjX35Bs88NQljiZ6nH9h09lVR6x+xNkYB98un/VnFt
ekWtckIIHD3z64ZIFXgik3g5fU1z/5GUBQyN94YiSfAXgaa8iGj8TkqJT3Aqsp6tepbFlzHWjYpb
+MUL96XgMu0e2Jpk9ecwdGCZ6sZTG/KMO6jkqb/GVYsWejyAE9lLcfS5SRHzftHY1KSx4nsRlQK+
ymz4soyQhVxuCEkn9pJWi9StOgrKJCLz3soLngpSruGKWJjBMZZbS9ottUqnq4G+gThmiU0EiLXE
umUASfeuTXzCO9TNIfkWpRt+FYVUSje0mJt7PhYrT9YubmHRp6K8Sw1v2Fi1E6x9qXt2zFePbvxg
ol4IRQAwqBVskwEn+XrNdBY9zOxiRczKeNni0sm6jWffdQOcKQK4o4KrP07ThO7fTi/ly0uZuQl6
jHcWmzHPAzUP+P3zICIaERUTJvBhAdFA10nAoV+Ah3jL3BMnU2r1zX9l9VGZ7E0iWg1C5CS9Ks44
r3O7sSRCCx8pIFMYUzoofukQ0wb3MVjNJ6j98+yr74PkGHXMxO+UpWxVh7p3OsZ5d9e8a1pNbtWb
pE4dntHfUh2uVwsfPjQIMT2oskeRvHKn7gVHmZic4t/vX13Q3+73Cr3MHFDLhXq3NFRn3EvRIR60
zGKgiIrOxs+WdtO6MQQaXrSf10DtaVUPYotGAzqe+XC8AtVCuCOnXg5gyMew9mmFVroO/Ld0Do8n
WgmnZPle0x9DHhS3K/BELZHJ2SwjeLdBnsEP2JHj1J4mEkc32/H2CNZI7q8XD17V4U3Nrzd4UvSH
tnZ8sXuWZ4S+O0bkJRRWlfBn9fV0eUH0phNZp07+MkPN2YwJ2UbG7/z7mLnITc3dajPT+8bBx45P
TR4QIPyez8qwQxcmRYOxBfpMniByM7fkGMYVoJ7TPgjoO/6M5rHslrY08MIb8umZX5CefyBDrf64
JbQ5FU7N5WAk3abIksKxd9mRMn9sJ5Zp0dX47UNGtq9AVTRxCHkrcYZCatZbu7Qjoh6Ws2y6jYCM
O2nYznTyy5HWcprUZ2CPj2Hc7nwLooOg8RAFClfoXGW3hREc/cDxsHLnPdygZjw77D16VWPnUu8f
Z92NuJT4quKZa0fDYMtmW2tAsqed407S7ZXgNSlhb46f8kb/tKuvm97GYTS9Y5lcMcrNLF7TP8iQ
Svl6RSSS96jKqH0gufherHUI8gzjVhpX4YsPIUYixrWQWbw8+nlWOcs/BQLYIRD1nstfi7WKhbBW
5yBPJsvTZri65+VAthkFF4Ee5n6p8z1UCTfXAgqegESuNFUsgRtLHc/ZYOHEoYSMyw+Q9Dy3QfDR
1B44G8eh5q+9uaOe0rPTGKCtH/PCHohccNAF5oQ29hrYiMmK04dOxcxy9SLfaxnBjw+OWsQHVrXQ
lvmlcE0Tp4AHdhETnI0dIMxOUXTqFrZWNz4Ue3vgarbIJ4etri7L2cUXTo5ATVexklbuXUxFKUQq
SqUT+eSQuVXB4jSOL9PVEdjpXtIdYaUdCB/VnGHKj29nwe8Wiv7WTA9h4s0xfwf7zKcf7HELZnYI
Pwecbbbr6neU+cHjvNejCZIr1/lV40avyCCD8xyZkJTENpzoWRv2uQTDZuESDWkoESXKh6SMH82T
WRUXiO14mmTcGsxoV+CadGwbYdTThaXCUH4ZQsFAOHm++YSbr2GpJezIogRnXadtUi18W8+VbmyV
Y8wFhuiK7fYSjT4HRbtr0m1XXuXNgxNK2Rd87Fprk+PCKWxCT0iYm3Fz5u2Z/DV5VsgXYOEUoMT4
RGBQUuua2AwEp6Og3nWsCECMiBomxIEVuP9pIxys/p4QSYGBHza9zlT1RP2kXaXmotRXkJskB5H/
cZuSRmRzCKHh5egqeJR1gNCqc/eq8dQvfO/9NHLmHP5KNaQ6f6GFjOZSWM7e6TSoDbU1GgwK6XhF
iSS13+ScZ3e7UbrPDcYIQzoMRje/EvUGyEt2u/Gc5of4OYVu15JaJKo+xPUyxlpfwMimRmj0BqV+
dhRgPygRxCCIrmH9//ax62DDQ+tVTeIPq+my3E/jNzWt6jYlN8NZBdVOaOApPXB3bNfj8LCr+djn
lUR0HzKtkCLeJ705B9F9fXfwo4o99GgfCIq8D/j4cgYAiw3jN3Lv3WBlD54ks3ovm1bIl683j1gB
/45WcIAHYYn7uK52PO9q4ySiirvfdTnMMtap1PINowj2u3OZ7MdbAXBn6CL7KwHzaQjP8kJkzKLF
87ggCN41f2yVdJeedHrp6RoTwjWRhXgtldDYJz9baEzp2jxXzVPXdhQ9uLZnXVvNONmFaCE39zLI
c717+24CcclTDHlG5Dj1TY8pzNRVOKueZq9tKq9TVpk78zrIRFvQxJcBApleqJpNLbik+jX7Uo9l
d+7/0DQ8K71FPoiQoo5QsocOML52N/qYUkIr1+6LsrQw6om+ayxD2zOKeQShlcJzZ35Hwo2+cRd0
hYwGmH9XuuNtSaOfTb3kHrCQQw21786KXHcGnGa/wOhRBWUXj1TsYp7R0zQcEniIUmz0tr4UMlaf
bnf7AUiMyYjEwPaFHo3mtIpmAAI4Bx2BhbhK+++HSDMXdMxdGee34W+NzK9FG/txFTdHezQEahHT
O4yK7AQUvvUfbpify8BdFw21EpZCgEppF4ILMEMNzHg/BcVql/MF8vWq8h05V2j0E6JMQrYi1uWl
CyyH9l1oQ2nmS+KBkQMfEqeQIPqq9roknXydbhW0BvT6FbRDJJP9yZyVxdWI6zFn5GbwZW8euWJ2
Yfz05zHX+0aJMhYO7GtnLjK7K5q0+sDVctwCwuraTz8VIWNvo9h5bA1cId2gfHQZh4ZnjriFW7p3
jrTurBNse0GUueei9LwEBYMY/rIjfdIwSboHP/trIM4eQYGqJEfEHy401dGRwHBwLp0aHupVdGiX
asbta2e8K/XU4f7yvPbZXtaIEcvYmWcd59me72XJeEDEsXPn+3uCnybFvqCVMD+FzuoNx/K5Kp2W
9BVwosyvCxq8pQEmad5NmwIdfFH0IjA+lA6lb5Q+JLMGe+/kvSX0l7KcvjpIl8afbp65tGL+819F
n5iDtK2JCK+z+Pdx4jjlbxECoD3vv+scsHm1eZa63tlazlQ0kPCVPszGdsK3zLhHjiPfS8TJalcj
vnx4Qeg1qdbVhxpvyRLIdVc/KgvnsdDjmovgLgD+wMJRR35konmCTzYrn9vXkj/p5KEpNdqfvglP
XUudxa4MemQjUrsVtLCouTjKQhWpVdXHh/9gtZrWjnZvp82NNDEnCpC4Pvbau3G9dW+N4Lqxh+Tp
2rrHv8nxtWqy0xOjp8GEhNYUejDcKhCj4dg5z5XxbzgKtifN+IC2Kvoj3YO65IGEh9CD/wlQsqds
wxzK62MhZ6Jri34mdMxtiVFBJiLsryivLwBBEgtJgNl705o5siNBgwoYAoZpZU5+e8rOZsbKFgx0
Tne9phAtrkxfzlctOVVj5wLhLtk93JIkSILknz1qlU0qbLh0i4vb4KCpsu7uQfkATb1YmsxveuMe
AzQr/eQna/BCLHyQuQ+PrKWrzcSFI4lIj3e2xbi/khBM9g6fbHC9ntASMewWZgxYW3fTtNdsHXOE
Z6ipj2LJO3BlNzSm22DPdM2CDSpwcX9ElE7rZyGkHVtJeMPs5lbwzGXVrqELiQjkUyvC/y8/dZek
uAwR+gSUng6IR57T+OjBy6/bLPKNYctZZUr4XLozWYlkjVCsc+iL4+Rj6q+OUciSkfYhn+t2Es8N
DSgaIMby7XfFv8I4lt6Bs/eLBiuUtHeAE3RYFuMOgkj13U0zlBxohprAh5+ftqYLI1MHqhjJsap2
5kZ8FfFHuli5bJU+wYb83yHVWsN0TrAnWksP2SEoFe6y2dCZCpy9md6pb5cq/5R2EuDtJ8Vm/MrC
UZZfE8VsK3Pyifjz7A6EZV69iJV1Q/aKIdxzMQd677WJvDkrnNYK9qs6sB9GnbsuAzW3daE/JPCd
lECnZs/CpmW+2qx1UPYAiB2cHXZB0Vita5mGy10CDIddXI9Lj4RBRCFN9bTnzUwIFfEcsYEChD2J
Du3kbZPLKfANpGwBIpCFUxFDqoAf3vN7W2oHnkdVyCJpzwWHIsuOkLFvuSd0y3fjHpeCglLNtRtJ
NwkdyW8SODTXe4SUXgDTRwSoMTJyAaqXrXL4c/S1mRGvbmQl+jGVXPYhGrsD7wKdozI+Z4ummX+z
3LjSXEWPniMjOcQ260hPgLKaz4c/9gKfcSJVJJyiATb7IazAA4Y0NwNzVtw5J6n29oK2j8p67nbq
8C8eN4V3FlfOqY/Mn9u2D/iZ+WRlYKLFdFoqo8hfViDfM4XEg2jKxTsHit2OEl7Ojoz01/g6BE+H
tNL8hBhdwHQZaqKKZNxmi+1NNeo6aMftEOoZiAFwSHlNCapHJRBZWIXZqLiC1/hup+ZI+TLfhyYY
blqs2bBIWRQBjQ1wGKB3hWZ6YB9vAmF/QIm9JYUF4und2UHv4sTqgh6obTSdX7gCWlPbwVm9lGL1
WASQF9pq8BoKZn7/hd+bJ8qsUtGkw191t5n/XT+hOm7pxh5Tp87dSBET5AUPq3y6icf2maCcLLHg
kl1fRNtnIN08hKlTPLgi/sicp4uxVxt3IuWE5bTHtg8C6U+E3kU4cvxuOP1OmQyHlhZyedUQA0bp
V78vyAmQ0dKPm0yaKgNmInkmgZ2FiYVVc8/kl7To5s1aQ5AwZ9htwjK+HcyGjfS7iIep7TT0dK/Q
4ZnBLwXkD4c8peSa6zYceKZtgyDEURExnNhMtLBMAXN/EyDCzeUk1Sej2ouY2ltkC7kwX0KBO1au
Xk+6s9bhbj4UJq/zaHO2jE8qpZPYd/NKWVPSkHJ9eQxoX+oLje9I7R367Ld2O0s5v9u6XfwaVZJo
pVt660llJTmN+pET823ryAirQCxsYOnpmWxn9CkC27y8Y3B6mQ1otADzl6hTBztdz7d0uKdbUA0X
4wBtV4QljsOaeLVEq2hx7Yl1BpckTPwXwfNw7HTXt8pJJq8219peB1fmMZE1MvzEnm8zTqzbpZvV
nyBaEGqpZl0netdV+GiOAcCIt4pIdk80YheAat3pUuhv7XkMv1umYbNT1jW2WsGAuSHpC682H95O
RJ94/IDM/AHkBBj79s12atZ/pPqfTcc+7D7CQmBsYKmFJsZXKS0JMMvNflIcpQKuzLJkV9Mkj0nv
haELEdUhy2q5fvhTE//mXu+zMKhJpu8uuaBvaMr/He7rkXd7zBWPwQzVDISDFpuv7Piwu03bMIK0
GDDekEPVv1PKO0PUtjYtmQkdHhjiwQlAbkt/TS8MpL3fk2n/yNcor6nryUijPIcXD1BmuC7Aaxxb
f32PlIO78QND5v9HA9P7662qhIySZ9FohrbWVF9ir57oUFGnqn7h/uOIv92m9xYIf0MIepniYoXy
qCirARPZKL4R5CA6AFjvstCg070fsGKc8hYLMtjKiXTlTc+v8CRL2sMRqJSntqAW0qRS7y3S22/Z
aYAr1LVBaHw3Ha9XJXox9w2fCqwi9D5lZp9tG0s9Q3pMakWLG3hUICAj4ggBa1Wz9CpISIwTiehG
CJxqxCqjPT8aamMQRoHfcZImIRKWrmEy9Ut1XEx4EsEkrGE/G17C31umz+Qe/gNCWyL8J42zmJDz
wVOuN9yD9mWMfQt10t/rCkgO839ysWOH6h4LWJc3rw+FhIGbrDL0u9dWeEKHsyvW7uY7GdgWLYU3
ff+AnL0E7WEvnShyXVReaWxkIYluSS9GCMQQT9Qa6sTnoMwKfx1C+B6mrMniybliox8yH7dAAhO3
WEmXrrF9KwjjIvPHfIxlyv2KFOsjFnH2vH7UhP7cjGeFVFQ/POO2Gml/5saDiOVt6rWG2dq6/uyt
wiYQvLU4GY1t4UD0Qo4eqBcEtIz97PM9cPT88H+gKQo+VN2F+3l2DLtf/Jsmg7GP4OrlpgVSgrZH
WzPcd+8c3p/3jJM1iae2WKUbI/uDfbHxjU6NpfrLaN/+x2bPNUJRaGxNeQKtuGeQ2mCrZcGjyVpV
2ScgBMsnWxHHkZfUyLfuMyIJS7fgIdP01bx+AqfbyL8acIMhl2Q7Uc84r6Tqla8Jea2Hi9ZdcBNX
mAOi54uIqlC39ParzMwVBmMXboHvsp6jIGkPsWIJ2BiYFTnyxqxa67u2/VNvaF4cWL3mQL+6dSMY
fRTGeaj56kl8J0qY4hFcEQwG6fMX5QLAhVp4rfvUaOr3+ZemhzvK1j0XPKFlLUYaWhC1098aR2t0
lb+mTMaFcDyF6IYmfUK31EHv2YF/DmkDjrYSqIua/tkKohX1HT1GT3QZfU7mXhPH/9ZUAKNY8f1M
jS552pL6ERHgsxF9Lw82ysA22LbXfcw52hDUmqy80QLOhOsJFvVMoYHflAH9wpbx1cY6wk0KVA/h
H97R0tnzigcElstuVThD3gchB67JlHcEoJDAqg9sWShBi+8Rjhay46mYAx6rCJus5MoW7x/Gd+ej
MZQ4WGHjGH8N8FRI1ZDoNWzOX/9Bjazeo+lMiyQLuqceljLz5w8xftRs4j1DKMcoO0rLhJNW0TXY
XPC1iR7r+rA7nreokiX0YfZZX5mLUYh+gZ+Cv34k/iqzY11gad7kh0EGktAiVdTKgKKGxccmqIeX
Ig+uVjtPlWjAyx8bByOS+FrgKUo4xif/+YawjG9y879kGZq42q3fuvcJcDO8xx0MtyCEYnvgLr6E
Y03rJNFfjli6iFZ8Bd8Xmy9dkz3LyoRdg7VZksM7tef6Pf8s14WyIWDzf4bU2D7HnXaJXAEliXKh
XIfKQhzkz+cEvYs6GfzYwPkWcezeEiCgO1dXVjeftJG8NQN1d/ZO4b3xooYzTfd2QRRiioKzl3YO
4elVzqiHJVCt282uBtLtO5ekYOyoVulWFs3y0fW3bXFFCYB14fUSGwRzFhXeuacW2swpILw8y1d/
mSlYj4xKg2LNCG9/ML3QZ5AFcz1Ngocuk6V5tTtQHrBZfKMsAiJHjIzRRsiPax7NNEYtJkYm0tJM
NRyxpOE2SbEdC9Zsk/HjXEobv9ZEKQVFBFq5Ifd3VONzx0GUFgWmCZLfMzkt3GSG0YS88fMLEvgl
4Bc/isewVZI3h3xGRik93WqkMKABMiBF7IATpqZx9MsLjGzsTwwrSUzem7HCy6dZXH7+0Ejt6d1s
uE24CSC8dv+hdgS82wxelPRtrtTVv4nWTUlNFRiTuiC1qKMF9g1+5O+xf7ukX9WLAAG3itAoDuhe
MGmDYxH0aouQOwaP/Ck1R77xkQRUoBBGCRWKESNs+KA/BpfgkmA124nuXFRxlGR2nZqayjuxN8ju
YbjtJjX3SUV5LyKdlq92ODxNF6wSuwANLWVcifPBrpw3aVDZFwmUfqs1ixq4y4gN39Jx2lRrbhCN
6jzg5hWZ8ECJPAV9iYMeaVyj0oLWx+njwJ+zanZOcoOFVnVp3NAJWZshnDIeNzcygwKJE3qjN658
8/n3kvbifK04YVVnioSbnXFDA4QHhYtOMZ2QnmYge+l4Z1nDYcOFgdRWgzxRTnTE6AMLcrnT19T5
ONgG0iRt9og/vk1iLrXOGpk+uVrfchLHbaLyG/+8NViLRb8kcXXhCWLKQigrW6WajSYB3qRT+lA+
tMEtL2gVdSczrqGsYuAlMN+7lqCkyweyi1r5vq+4lUOX1sLzn5zbAASO4xrBjqXBtjNbbPT/5co5
xUHlR9ukwd2YHhLb1QoYMRcWCwqeLZV7zlgkn4jUCWD4azaXmTDRfjcqqXCnXZbew8p26GEV/Jy3
+t9gdxMx3yTCROw3ktOB5tL5p/Obxjw2xPiKk/iNvXdBP2r3qqqq55bhUSw0tTCGjmHtoVq811vo
HNqjMuq+VUdP08Pvsxsazbt1u5/VXr6rnC9kjeGmYKiFEb9/x3Bv0jzgPKSJ1EEkQdtxzVRBp3C0
mHJARYnacWguabDN/JLwWe0SSrSVRPbftoqqazlfkb5s3wQI/JFM8Z4A76n7hI7B/uNZ+V2L3Wtw
gmJaQd3Rvga4kN/43io/8ZI39Pe+J/th/7wsfeI74G4H6FfJcUeqHwoEFK1J8LM8MWXGw/R9Fie7
DZPtTxTvdGA1lEBapcJz4WyG72IF6d0dydRv5BnjykeOoG+sElLqzdYkz6sH7z3FTqEfbTMjSR8C
9uNPfYOyY/s9aolNSY4fZYQO82HYxYVOKwkrsN1Y7F/w4RgAPaFfv/77ct9lzCF1xiCu5glFEPZD
368vxp0uEiKgkZAwSklKmVxE2aFH3JnwsjZqqv3pBNAXZbgXaqJLMhNv1+Ji2pHglpzk1xBT5ax8
UL+448io+x0mmswA6TK3Xd/DCsyVN4bs9gb0bgckMy8tQ2296KqujeHOAvGwm+C1HXo4eA1dUZ+4
cw6WSJJlxUW2Qp9YdbaToWj+rglOEkfnZsWeiqOfc1F8XXsJFKjX3HRzwrBkr0sQbowWwy9Jlq2v
fLgAsUKbiwgr5RphVazCkp3q4VuWcnJOn//DXi7JP7d2Tc8s3WNk/UUo8TPCDqXy4Kfv18qQAAbF
YVXfrVK3whUR/FuXJPpuYaU6X/sdMPic/a7I6KoIzlFNZDVO+oMSqaK8dhG5/GMfCuQ4HvoI0urb
qbr5JEweFc8xgAaTavGnWazvZXyxLle1AiOwJytjkxRPMSVIRl5eqPG1GXBGv62BJ4ZXx7hP/FTM
JINmY/QbtehrEY3gClASCTyQrtMNzxfRSxjwhECmjhqNUJXNGqyocW99xnVVZAljKHfFpHE7MDC0
WLRBWlfgOkAmGhhD1WNb03kGFOjnHyxrQPbj4RyEKa6CQDmC/171p4lxei6rIUIJpyxvC2q4KIa0
+fgnBwE7wpFMSpKK4nmgaM0cWEoe7M7+JY1s+5kChui5eFmtnjj7ZhMYEB3k1WQn9h4kSk7mkny+
uWDwA2sMpF9stpt2MShVuXaYvPq3PpWfllcv1rNRPrrdoteB27X53QN+SKqgbaTexwP4fqrHD4KA
bUWsf/FKZv7J4r5fO9rm5ELzv68PmpaYwipg/SWLykPzxWIhUTmHINFRNt+sLSKkqBLq7wXlORVS
/UqPojJSLo9Zsb9qKaNifVe+g1h1qm0GqFPhR30oUV2cJ1PuqtfRJ4i+Gazf233A3H2rGhSHHRM4
xTmSVwiRTdKOpR75dHtSfHjd3ylJpTrCuT1KCN2e+FF406W98xgN8mh04/5uHeofJ2FGP0xGk9qX
l4mZpFV2KmR4DiKdyv5br5f1RqA9SIMRT1bdCCtSoiAM3ZuSROjCU9t+hCGlEjLg+uP3LHSIWBPJ
qYAgIlMqKdR1n5M+gsVLCCJSlI9J79Q+OY0HcGRWxpGvcx9LrYIAb1MWJUzbHX/NHT7v44F4Ee4h
1a4pFSHQM0tJA5HIvmq+BBvY+gLV5METEyH4Sl61zT9QUCDRmtKniZK+SXOTJ0g2EaKWreZavg/X
k+5lJWtBkG8MqXebO82inZLTJRjPUBNqyxCYJFGogYY7Gqk5MutHoOdAiCqkJf/ZdgQKyU6lSM0m
Gs9/PSK7kBUnVJ/PqE/vsyL0nVMr81iJKyjawN7qAh4icn3nOc0AvZcD+dm0R7n1Vw2FoLvVxoGt
ustH4L/e9l/57zDGLjiOYqgxWSu57e9Tyo4QhCWqRR+Mri3+dCPc01k44FcuPep9z3e8sRnX8mLw
2onFwvlz4tgo1vwsN23mnzktA0wFI182So+7t74iHb5f0+k4Tu4EEj0iQJ5NZaejJTXYIZanuZdF
dVnoGrTive82vbzWV0wfB1vuldujoeTtqKslgOrJHuJTcsoTwoVYi/fM/rVUXoX4PyTdrlMzXCws
tA4beNCgDSGKXSrWI75P2foe0F3hCbD1+YQJfFEK1bcZix3bEWnJIUgYqvyLd1lNgZdvwFxlHUzy
IqpDz/sWE0vA+gmxLwFltorJHSjtNVTtSmoF31Ae9ZCPZhW/CPuUpoFo4tVqN66yEqJWc/SMsJpU
9EZAULNFh+j66GpNIbOE940by2dMnfj1wFXvHSX0ZQxDtivbgwx+VXEfvt21o0VZfLFCfTmyJ7PZ
dc1Q8JHalQWjuLei8kkZJlS7TcyZnLzLj844airtqPtyIXcIa32RBzlE9zLELaK++zm8oBptZLPI
GRYQx2LnM956UBL8YLcxLzE6K3dwUK+g3l08oQEMESWmyTzv0vVsl2KESQ/jeWAa5dwz6/XNnt4G
M6Vx6KXO8L8t6t9hFnOCGU9htIj1NzOUYo+U5DOcHwJyd25mt42DNtbq/fK/BG9n+8T1BdJfPxIz
bDU5PTDNiK0OXoOX/8HL8luKHdY2jcrEcNJLgtZd7b/5ivGv9C+LeOQ+l08Hbu7p4tFrIcbmsIKa
gJso0bek76j0ge08RU1+6KtymU5um/QNSBwJIDkpBbTOfTeSf8zzwgHHvJMdfeNht5h5/V/thy6y
8ua6jleLutjb3QQDdNCWP46r3N5JwCQVOFB4+bjcYwknuqEHPj3fi1kUUundafiAztdLKg5Q8jMa
8t4UkL7ePOx053DkHq8BSA30iMhw9cNI66EeII99n/kXx1SvIz28Zip18uTYiOJBjzwRgGmF9r8p
zjToz47w/uemCDfbr8nCu321Qmetje2p05EDEdX75qKkHvwzaXRwROVfKzGAJ/yU0zCfIUcbNruO
ZkH0OSLmxBtyIvpRadJWh5HGx5R+Y9ZEPvDNJdvirO3CxnAc4z5bvReee3WhH/VJBu4FgckuFb21
ElLlOhhgdHxXopAa+mzmzp5AAID/ET13TTWelCgWaCd7XQ9Z1g4nO4scPsZsOuaDpKoYIydMpB5I
db9EEYWLZiwy1LKZVtWPJ/+vRcFcf0J+JJlkLMQnJQgMvfs/wWLE3I1jSolMY8cg4bsUiyjhL5s2
bWuA+aH91VKD/cBPqK39ULR9yGaWrfR/giJl18w3Sd1KjGMrr/mV0JU7VsF/4eXNAcUl0Dyypw5g
UTIe2vpsX40r8XKIiBo9wszgt/NqeABBU+UPTv95HXXl5S4fiRjh7ozn7Tqez+q07OF4dYhfZTHY
lPcSwCbXaRPHO0FojtT4jH6/LuBeD57d3RU8cYmrWwqa2mGMHcIJ46UFZ5mE9JTA12QxdSDeKo4B
BSm8OpVQgQ/unnyyO+xPZi4scpJmSKrigQ5E15Vv64bayjOR4fWhKxEOkyT7sNWjxsidAwbHjMmQ
GZ/OnyDnMcS7LACx5/jOLDaCsvKtoaNfAoQGNUNZM94DyUobUSA3g7ArdA1+K3AUzRedb//VRLFB
3X4TIl2blMgfA2N7tr0albgr1ISeHgERRFbkTlPlqkIx2Ovdf/CQ3ngC8RM380iCBuKjI83IAJq2
5NdoLLXmrAgXWfbOhBSl9AX0Tr54WB69UTg5frXNvedw80FjXyxx8jvqUAVVoHqJUx9IhoZB2vbR
OUpcUYi095dbSyyciiHQCAASaEczLCnmg7zjIcV1UwhXFe7u2C3KFookgbEf5GDyUsjJ8wLdM0ty
jxMLphRmdT1m8DTJfV583NO46Nn86ko/wk4Ro+JCjJZSOqmv0rGIocut4L/3FJPbRO2bC1xhRZPl
QaqF9Q8dr8aNPdPAk2gmRKMR/grZnK/9agMZXoZCj1HTRUGRItpgOpYBL98SwAF8BHNw9pH7sv66
nHwXalDy/7TEAR99cFtdxOshqKWeY9wKbzbGYCkx1N8AjYfK7JhItT8pQ2XartZBeqRnuRQSxpKF
FZDM58kQN9fM6Ar0kQqLrvfnx8Gz5zeGBowNh3l641iGPnIKSp8SN6v3dlvlWfVrH2+lTyuWP4Jh
qoxyXfiZKz0WW2NmkhJ6txSnwVTSmXAeJnoq9UHUWbv0PU2YclOpx60WM5DZAaNZ3ptTCYmdiylp
FOSPrsGU4RICjwCmXfSYYAg3NyOrHJEP6hM6Ygub/c/8RDpyo0DtgBcQZLCV97MymQheTpkhFf2w
8vswfnNiNeI2BNIM727kvdY/s69XOo51GqAsXHo/UyHdVbs0IHkhkhvWIydipQMB2DC1YBN790H5
zcLnGzzdG+gw7B/NXStRs8Lz6VRMKsYPkTJb5zsS80E3PHCMmghCtDGE7mCZEaxMVQI2HyH2nGrf
HjF5QCXJMSYKCDaOQkRFMAnkTsfSdXdX7avjSsSafsUHw+664CIclkIfiapEQdpqfVxQQdhVSWiz
LIT5t/dhh89ZcBjfziSA9rINcfbfeDlm8SAdhrKPMyInOEltS7VF94vVDc8zbTBCyXzTBhdxLQyC
49rtHjvIDBqgBEmmoAGrVCitrLMLs+04fzKPEEz2pYAKXz5SXz92I6blVoS+dXArGxVD62XmPorr
Yp1kr4+iIZ6b2YBUNPuzaCJdTFDhFXtPEYywkI69lrCCJsypDwkbdoK++kJI8w1gXvnqx82ygFBl
hlD1BJ8tMQacI+25t914SpMuCGlPtQRTrbAxtRh+VJMECi96xhu8XlNQQdYjkcGYMt+HXbvh6XsA
NdLYMFzD5Oxqxp6irePKLhsR/ijFOre74RJ7x0I7ueCJIdQUYk7L9Xm7xQDxqnKJzGNr+m0/KZD0
nN/4+XCDHL2UTPBLBPfEIyQxWUQnBUkvZHeLRmyRD96NA+mqDe9QEb70NsDxOwCEZmrZGXya57DW
iNIdpuhkqP8GmFI+31M035IdhV14NOe7Az//NVJSDyMT1aFxlk3OtwTttU0E4zM+PdtJPsHxVI3w
gTHkWLr76/2GLsMW7vX7VbOWLRbplZv6yqtemsHphduEewpqgTKdZJ9Zb+N8r0NxuFYBgFbklePI
kjdcSQnYaFzbgSVPA59z4pZhz7ZbrUsHJ9DcW+CSqgGzN+D5md1I2+BRn8gCUNUtHjkmPG7odBdF
7p6BYNfEfILrbF2/g2IqYEgyUywii82B6c1MeTiQk9g8YaWW/dm9/hO6+NENjYyeZMkwt9JBLVHR
ZU95z1FzgTQYV6ugPKFhrOx03gD+aAJoOw/RH5N7KSd7vP+VMtoVbMEHBIp+TBlgxOxD05HdbbgS
HsZckeIQSC3Ow2JThiYlTpkYls9Ngl50YZOanV4mDOJVvyUeMe2biIXr9ES6/AgTaYB3YdNfN7U8
J6H2yTpXdsnP1xPV/QcNuVvd560eZe/+vK2H9UO5w7MuGg3j4ImFj1c3PC3FGB0GiwgVcqEwl5Km
KboEqKRhKdgyDaPOpuJ3pC+hizhOg/ydS5f4u/1qDWGWBUw7y/h1IV/cfyyBibwR3NZnXvijnJ5w
UnMbEfRh0diMKHHvvBrxNScJBre1gsM0eqSB2QaumKF10UCxnZQqPB7GYu/1ixMrpfo69+XW+izx
NPvJ7iN05EGbEIvYmve8tgSHT3zcpvaIebSEErTtJ/zKib14gtBho2fhwg1v4U6urUMzcKYeVROQ
sSbOyriNcegr5ZoW0oJ4Kz2AvkZeiIHhhv8YGAPPCGJFp66U2fnoiGuk8uGPSpIZQ+RvBTXcbe1/
1KyoYE9wJcgr2nOhEtLphO8RUkBJAs11+wZrX+psNXAU7OV5QTNOa4llH5asTuIk4ql/vYgRlw2m
7JuOjmzRMaB5hmgT0q7wuckjpVzm6eyjlEDjaqMhx2PLUZm7il8hebH9jaEfInKYe22zQqR9K2s4
5WB61dyCTwEATf8AV75QWzIEZ0b+q8+bsRIcqrEgJu69ka0CTtoZn9yPCxXwexSBnPoAms2Z9oKT
gxdKanCOUn8ZUHvWzuoEb76o4huVabbuGuRAsecN6p7XZMajx8O3S5fxWp+LdccufKMpdbeX/Z/w
4cQem4DyuLgWKuZalI9tlN0Mnky+KRqCu7qJFDm30nFZzPPMtEMqaUgNtYxSRGybFOpCVXRlTpdg
tfUNwOW7JcRpPa6Y1ZzlnbrvMe2JaJdll/gi8yBS+bLP9cXMcgKYC4zDnn+qRZp+Gw+lHdjn2Koy
dTUDsFxpxr9g/p7DB3aVApt5UjlZ8dE9l2v3b+irdlSBU2ZdTjRtJ7LcJoAlVZFrmBAJ4JeWuNPc
jIpTAjT7l8WpcAwm78pwbl3GqEYZvQLMPNZq/B0qOD8iSoKkGN9Q+5VwL6L1+q2gQd1peAIdafg2
F2jpTjylue+lNLgeMcrhoR1PPDKILokZW0V1/CJmz0USb/+zx+VgmlvGtfp0sqyLiwsqy6FiBgKh
LwL/h/54NJyF7KWwaEqXPiJI/cJ4v/GjAU9aiOnKsTIq9MzNhERuEg4cIY+i0Dm3g7p3RFLPyfZw
4OBzwvN3sBame4Fiqc4H3nybLv1yn7SY3R1LuZKRumIj2BHKxPCmc5+ScpAAQXrWFjV80zTw4XRI
Bv9xZBuTpnY+uq9ehJuV3t4cVltNERJ8wdK8EPa9jwvVx7fSCumlAstQCvDdGG3ZHKtyISGTbdy/
OgPzxJbOeKfjApsE4mkOwewaJhSDg7cq3B7ZV6sXvOwuJnayZXPOCNYCzt06c/BKMQOHUVQ9MBTu
2tZLZEJItaCTERP/vilkJixGWRQqPwMIpvNfbGAlqoWF8/uYsxu2O7dTUddET8xgsz0+7dyYQzfP
NJhe/2Bw01pn5VkleI6EXQr6R2oa8vXdmh2N/hnNbksVUtH4BEULSu2VpHR0ueaHc0eruOy/Gu3T
3WiLDfnG4YSXVHeoHTZNdGnHClqZJhPX7Kmun/4C10PKEw57rFuB5Fg01jceT6fBJd6LVPBdCTrv
qxzRdNDTRIODmalWVoFnS8W2BqgAwTljKqnsX+b0dHmd/9FFLtflWQCBA3zE2Crq5LvSuaVmPpfF
8Qs8KBmFoEhXyiWO2UKWxQlg+cD9RBJ8JCJLaX8DrFB0kzY2FS5RKUhtcwd555B4tKbUgsR3ug8M
bCFVbOlKcvRBcqVkuUAqQ4JCDhWeaNUQ2wq0lzAWGQt3wjvKB8Ke1Xaid6Z8ImRt9ppXrJnfWY7M
WJBCgW7w49XBM6xZTeumIywsMrFueOGepDtWWckdCa2Hem9QvFRYavqc1ayLiSIUe1KMY7VqPJq+
MWqBCElBZ2b/kmIujlkyNR0k/610p3eA6ZtGNFzjym1XlBAY1ZBRQlcYzD0qy2pGkZ5ruGPcKEd3
TmR3Umwzs5ruNg0rDXauitQRj7hFoRALtkkPBtzHjf/Dlvkrc76QskYfpy3U75z4oxND/gAI+4JL
6RiS0klXWxK88NdeaE+MYZlxG61/8Ut57XVsX4O2QwtszRJysuVaOCoNLDFrFozdNFYRCn08n5++
ilqVfbGMcV7110/fC2EOYGa6RRzPmNA7nRQiaUOlOc4g0lgWL38QnVhZdIjhGkuBC9XXIhLgJMci
eEXiKjg9k/W0HDlp1tLkrxG+bB2LiHK3a5J/qQK9+YkwEPpeSnT5C4ZVL9P2ccAFDa7RKIou+9Qp
Xtv2w3YR5/WWljLTjubq7rAs6xy9NY1VBpJ7sWuWL9Fwl/GD/DSsnkUnev4Usr+enTDxlx1Medt4
rer3rmF3BIGtym1/2l66ZR3munp+NfWaOVQnrpuYiIFrnsNyI6YNMnYhHygxPyUGIWW3AfQ4ePFZ
nqAwZaSIV3n1+g0xGoHal/j84Ku5tv+KuYUiJ3AkERfoVb4sMlI+z1+Bdoeov+65DEQhXfgubaXz
ZosLcHftlRd5IUZG4jSRWFpyFusw+A17qrXmE+hLVpCYcnhV8FI7+Qm9BUgWNZdv4ZwweMXOaItw
7ELwe7cywY7zV/tGqkOlRxnIcb21KzB/vGrjNyE5h5E7zUOFyL4A00/GcznR9Mlr9rJ7mQzdOSoz
kX2Kr0glki/MutJsciQPekQH9IaCoA3eD3L/XuUE2+JcX9tU/DPMsBM0nCSeKgWIeeP9Aub/mdA8
yH/PE5eWADrmqJrt+Gl7dNj9rnbhGoLv1pEgggWvR6KBAafNaH+RyqtA02bjRj/2mZvJT8jQ3sme
ahkHaedcOUnZ+fwq/ngHKzezF4Teh4PWwwCtuernFyexGu7NXCXINoy/ri7rMG6yNUExEQaH2PZE
MbZEvm2djYe2Uzt97Pzqegqar3lc9/E3+yncHuwuEa5ZLnsIjCH/ayfV2Gd7L55VhBO8ILbkqtmP
433iGksdly7UFAvpO02EOs3kSj8zl+N64ktDMTLrK22WuUh21xh0eFVV8H4LCzC2gULPNicedLZT
iFaf83YneDPTx0X+yTPzMo9ITImKFOTIrrQ5Jec9GmsJh404DEZmW2HL+5GaCDZ3UlDz7udyvmCi
oS8FhdcCCmMGj4o6MBmB6bLFquHBZY89H321OlgQ/udp6WHH/rQLrlTuRupBigSvENZo8LriSsvQ
nX7huLeGidnpnJv5sXEbjOGdwA6OVu9Ufdgii3eSD2fefktatyIDSg56f+Qbh1A6Ee35RhQY683B
SApB8yWpx01tZXBjtsDX6X21/oNCG68segoj/0V5aoKpGy5TX3L7WVjeYPC34k6jf3zeTc7GjfVn
sGRM7lv28N5mxDcYBf/ppDOV/5WWBFThw8GapNPneFQCMpqdIM0R43/QpVqmnXdfV8Rlc7IX8+gZ
9VB3t4C4f5Uu6j87IprobNSnes/+NmSCAIJ/fPZKFk+S/U+t+jAwSpDAiW8bMROtLHa4FeiHKesp
GBNQQhtvG5XrJc4dBb2oJ1ORN1fnt79DxM21ZPBREclYV9+UR/hqCCSW7S9gg+ioe/Dm93rGLyOn
rEFYuuChyE/tVuuS0FcYcb4emaMzjG2DNGa+MM2TwDANuNstE9m3bFWIZ+9tuyVVMgdxn92g8ZEI
n/NAJtySyU5wIR+bEfsePmBxN/xyHcJM42EJMV89sUMVtnHpyGBYdjdcSi47I0E8kTITjyvNqNvu
7McCOqQB1xfMrSV+xj0D3l6HCmp3sDH3Siidu3EiB0oKn032fqcEnbOOhHUcfYcTCfsaHbHIwnrx
6K3z89NWwE85dpOC00H7CP/18AuzIJW04NWK8cva6XydZb/7r1OV3yjAJjz+t6PDbs57+5cYtSAK
eiwsIrhqjbJMoTt2RZROcNQWGM+UZshmbEr0VyTQcY2zQsF+ZcExVqcRtQcwT7XeYDWD3ebkuQxq
CBZacOtfUjNtrxw3XG68HmGVKL+NFQfeKgBEMH1B7bck43DG+tm2+G5cvs/6YhLJ24YMYBgSmKXQ
wxhiRbyqArgFjvIY1EF0gWy6QERxenGD4wxMI7xGRfgtoQOaPY+6XQofaz3iaa1opv08U5Dl8Y23
37f//CsO6AnkjPpRPKqnynG39iD4Vl0Ho6BSnkWq3HlEbBrXZvVk73UkVdzuhPoX1qTJfCNrVH8Q
sVfg9EpABIvevEM9tGAPdbFpURgKJmSh0E+nrN+2EJmu0MruSlsYl127LmlO1AAjjJmE3XMjg2s7
up3qYZsArSclWZ0CwGzV+id0PMxOrsDgHuqJ74ToXtlw4gmMEqE6jF3WSm2Vfwp3JE7uosEaMM0t
fqHnzVDsgdDzsgWmHZUf5EToB4I2nnEd2Msj4NVq9eJxkj5d6UFzc0th6aKg4NFr5n4jInoPOSqM
tq7iBoFC+0GchcIs+BWZOm1swVt7W2g5H3A8uqecQsrgZfFVhzKRsHDJHfPLnPOvR2oAF+xndeXB
6CvM3Xb7/DR+2bhsiI7T/VLXRQM45pZw5j7jySJV6p1u/aoFzDIU/22eJlcmcwEV3pFIAjZokkIc
T5aVKD8DLp3hNt2Yg5js7wxP1onfdSgqQum2N4WKmXzNxtvCWG+hCNQAIJehykKfHRy4DoCo60vD
wJ75HkQ9Zw1LwHBiz6HEuMKT26Taf9pxBT0mMqboCN8+lQrhc14dBFf91/tJMw5FgFgWVIyXFw2y
eC7Th+es9kRUCqw/VS9wAzNdj3ZtfF5V/RjcoPUv+iKmpnHTHk6cRj2QTGDEwpZ30KG7KBntsQgU
e7clE7x1HMaX0nFniOj8X9PgRIE5RKfUq39HdlVAYwdT6H2uGMes5mTlqVDDK3h+t/lL/DYqG6AY
RU60x2Z5LrlYNOB+rbhOa3cL9hn0gXO/qWlPmbvXZom91Z4DAaNdQT23vqPdzRn+DASEKtiqbzoU
i4HdQuyh/LeueIlzFHT8tyKPgCoRZWwJu7SaALUqiWX+1xtZcD64qD03b0xxiBanHHTU5F/8M2s8
ypu54c7j3sushez1GgT8wtEe+VpyAdubzzdapLEB3JX2L/kNtzVh2to3y/3UEeBBgCdh+AVGE/eO
+keOmrDdRiHQfWH76ihLbs91yrkbTag1soWBmZmFqNX5IXtDkA0Ka8EWmxVTe/bdzOhgvnUwPptn
EwnqYMO+aEsncRa30JyNBY5M0wE7SF94HxHUwapJHyIL7ZdrOV9DScvXfbHpSxYEq4cyvhtzEM6Y
ambK3bRTOB1OPSLdlCNzefPd5zjZrVyzEbZsdwyM5GfFdUmkyloSYM1SsttK6ADL1T6APLNCF7ZF
HxBpxBnV6DplZ5LicKLeSOi6+rihqdSZ3JTU0kCYqsnrMgbHyj7YKJzo/kM6NQrJj7Iaa3oZTsH8
D1u4KpEfLVkUCZJ+eHjw79It1sepx9kUCTMde6G1gMAlf8RRyPR7YIWlqmaOHRdy2uRRkyGJHFCn
wS7iRe1knUxiWRnLlCPqcPzFglgjn4SDB7+9Kc1Qkm06ihvq80WbdxTk6oJDCTVdy3eOPS9VTfmz
WdULwBH89i8NnTLojl7sdEoVc+WcBwXGS7HfZKSahpdmwYlt2hpetVMQz4JTOBWfm6hS08SmuyvZ
qwvAuB88R9ScAUVrRji2T+HwxNN4TQGQfU2wpa7AcDwiikJe+SV04ryMiFOh+ILbfPwAO3geKs3H
t0pG0SP8xUNbKGFuPzefqIfD9u8vCsyDJjQvBLlCRXY+G3pNvLM18MU4buEMfD5XOLxUBMAox+jJ
+O3LPE/kw5WGZu5UlAnuwy1U3nYQqac/vlFrUaPv4spWa/8LsWBwI3J94nzL9uhlrWx/so1OPOvd
h7q7pAVKRnCop9qsD8whqdd+Z/IkRHAtrNNSekw5HgSMHqQJ93tUt5nX8tKOOEJIjEKdcnWwfUFS
CiwWUsHncjfIZ/W+Hmaw/ybjozV0Rbg531DSSClqwJAtZT+LA8/5q8QWq6guQP6m1BaajcvI5duG
3iW+KUPjHbPMWsuJrv8QM4hmAhryZ34qngweHxtW0MmpPc+JEwNnxp0+9G0tBRXLAN8BRdbtzd1m
Q/vyri9+iVjdBI9rNlo5kVg7t3Egsa3emag8P6UhYwt/scCYb4Ml+3kttNG1c49KDcWKzWXa6/1k
B2jCeMYSSLjv+KfeqMJrk59oTXBP9ZnYjoSId+Ie7ND8KGLSZAkP4sc2Ln4O6wHU1CSjxHVdzKd/
63VSxIRW/di0PwjOcBfMQMFTD2nDAM+H1Me94fkG6+pWz20P/no6DNKrx8/swOPF3XeTKAIQuuwQ
V31zcjet28c9asOPo6ayFqisPK8cOWp7TPIVQslD5Tizc943Ul9IhdyU+t047EtAgapgcQ4TzQDT
61lMCW8DSAvyxv0ytjC37IDX1B9c2KC/j1cb0KJZUT5biW5v/JSHK+ofj5QVonlm85twxQlt2qWw
e8ud8dw69PxBFsGA6RrxeY3ElE3PKE+MA4clY0zHxQkcB+/VL9Mi+fCtN4RNpDz5UU09gEQZP/3Z
5Q7wD8fzw9XNdLuTmEL4d7AFKVY6TzuBJRyn+gZ7ZFM5PKPvvLXyYYjSpHoIsPrXBl6k57gU/23g
5DPr203iPcpeYxjmGpaIwtJbtHTFP250ThKgfPq+FLgqZG0yW/QVK3nYeWvuYaY9Qj8Thz0P769e
41C0Si1/jDjl4+u+swTVacAUwKPwWzECqgNVC74SHfE1s5Mgg149Ag2B2CHRw5sfQmS3WISaIoRk
J424rBp9qpFUs7z3F4f65z0dI5Hwm2YfHa5DUbsbuIDuRUoO5sZhS1GJgkOINl2RXCSnYK1JBm/d
cRwT3noBKginYd5RMCuOh5ZkMj/vobDwK+lE2Eap07LkQPi/jA5YG4fqtPGpN8UnqBfhXH2rK/G8
V6LJBCmLrr6P9CW0Ywp1iKNDDVqGH2caQElVBlMrA3u4SISQhAxN4onO2B7dSyBtpAIITPzRIV/f
6seFuKFpKCAijr+wktZVtICDLGHHVhO7vGVck3FBdHK+Mn02OmcJu+x+lZWVgEHr421acTTmHrmJ
5xUhtqV1jKMyq0jKxSkZ3r0yBeyV+ZXloEanSQUCbllOLdQdEFW91EMKRPh5bAnysknT83srtfsj
KT4gH7RZo9PDclJiEMkdntk7TmgsbpojgzEH/WlL/n8hCN8ROPlnO1Sh1DLOU/458tqGxHUEvj9h
CdfVqE/rYzKuAXtdidW+MPoMiXyxxO8QVdtEmimuBJ1xZiyv6PRk9cXZwlsfjRhUd/sFVs6jKrGU
SC/zSLMIkZs74GNPgdxouLHRqeiFy54EsIC2ITDN+eTFBpaE0qtUq8pZVqTV90jiOEsBI4B+tJQa
1FYqyiQ6eWlNsbZIN2qJsIcI8CDjQPItlE/8byukwvVJskPUren8FnfmIgCi1btOuFHU8/RS9xB5
zBh2oZlAu2q3OsS0QwVkJxVJ49pnah1abqQ99rcRj4HQKoeZHRpbfa4WDkKnORURsR1wTZlriwvp
q1wMp88vCF8Y1z65BfzLvO3dUrnxu3p2A8BclRQEmAHt3wwxBGu2wZOUBQO2dXPosVkEJrDmbrBm
EcyaC/U79JdmwlCBIk7xnGwVnr8joRdw8KDoqyxAl0E4erle1rW9KSiY6wDQIpfhTSPvp2Jh3rWu
4o5evMNkQmo4fvJaB1L93f3vPBNPR1VH7LupLijWrWtKaT16GDcrjeTNZS7gxAHCE8rUdTkZlYVf
Q0K2LbsJ8vLbGp8A01+pw5FgHb3mhUXQHnTIDSF/ArewNuyhIUHaRVqk4vjVWNbeWs6YckoohcOD
h1oBajHXUEcYIRqyHKyKWRNQW7t/tsziTdwGsgApK6zcP1q8it3Ggnk34L5s3HI1BY32vCqsEkhv
71KhheA7SlqdUouM1OP08aNlgqM/oX+oBDEfZSQjX88Q2WbEKOF0iWcbaLUO3Zlh5RJBiwDEu9b+
gyrER8V+Ezx8YMIXDOlBlqP7ZPemTA50HqkCVMrohhkwjNxb//Ijt0rOM172oeH9FKOTmPwK8xb7
yFq5fVtnipricEPEebtgfF/Jq/1LJSB1XK/v82MqemQoqH1XbM/0ZWxP2zXyF4lII9U8U4/17vsw
P62lIcGcBp9QjY5SsKRWPM8L269JIiuByIwowIitvRyG8hoLCezSQdzQYJ/eMMRFqheAKwDTnA1+
Kga4TE6TH+zw3bUIdr3nX38OieAxaTIE3oUJr7cMAppNVLeG3XjcuXqMjwJpcLmS6y2LMrbXQAUO
BvRbqqtmcb/iONxTqj7YWLRO1UL78fKiwap32UPjfh8bsBjdNDbIR6X5oEn7gRSTa870v/H1jVCx
2JqDWBDrga1UV0YqtkK/KR7m1cv3YT+DQkE11PEN4ViUicTozXEw8UOgfOz6uEacRrRDtzdEi0UZ
+pFnkrpww9KtDaChGMP+6S/fLYf7aMUJPwLgAkQNPJrbFaQEHowL/rjie42ou0mAZ8VnCdd0jKTt
DjylEl765miW82vZffMhI7lMgFSis7DfwVSHmxWBsBSnuRs7Hu7Y5CoMuYOFoZBT3+M61lVINmEg
xk2j4ypCDNfhDD3P7W1f+L+c9YRkpgt+z7y57ora2krwDxszA1vTXgm+pjB/aXF8E6QqRjcgUOeP
Jq+v/em4KFqZ2TA1TbcGKr+jFodE7C7Mcv3z4Xp+Cne/q9cCYCT2IXVJyB+FCZ2n99piUbktVhrJ
xZQJq4ULXiqQe5YJdjp3E7KYDpflm2D5FS75rR7xOwZBgfgGpNM/EJVig7EFAhMHDFKMVRo4bml2
xDui2T5XSUq7Yn9tSUGeCh1CvLepLtz3m7f6tVxN42Nm/U00KRftvlVlE/nkD3mklnNRCAwMWNfx
W0WrXdHlae+yNYfiT5yGKGl9mFSuujjeHs6yB4emqm+qCFUA7iSwFwApkChHtD4zvpTED2oBXZwE
T0o7AG/YzNNw4uperGR8fuQe2F7ct0N9e7lAZLAcuiaUJBFMxOmxvpbsy651iCcAawswU6Ks9WCc
Lp7Nk2Xt8Jwx/0sVojI24wuIORf5nV0zFLUnHm//dQrmv2Ca1qq9Qph+fj4caeDUqZqGpTC8/jsr
6Lw4iTfuY+YobA7D6WSssDt+IEVVw2CKnAfgZZpb9DIeZxN+7FghloRI0EWepDFIhTDCO5n5/bDX
OyVQXLrYwJy1wKRdr+rIJiJ1wIsmx8idE5wJAWpqVFY1+MryUlJFVOd82Zw19BavnwUAu9ajLkq+
xjQEgYNwKLg6iHT4AYBa6aZtztGazHawG802VVDYQmt5qbnbQpIYaFe6oLwLa2PhPq/sHBSsf9pp
vceszsJFFRdD9UantC13llMhpxnVgkbr5ZbdUpDEVwuJh2h/AdymyhmBD5YftTg9RfW4+apZJ2AM
RhSYOSOMWwhSMtfY0eIhzMZzdZOCrdt1JSDKyEKOU7xvTfir7hogh9VYicqX3jdD4GSLT1zguVx2
L6YWwanzXjRv2B8io0f03QDdvuD6ihg4R0S0Tawx5iAdVDc7d9vqB+SJGlWQSjZgGAN/PPtQnWOJ
L3MJyYCT14RsovQpuzSJCN1UE4DrIeU8poCZRHHhJeQZ2lGKlyWD/KVXlp/mCLCt3J74PiVvKmAv
IhO00ZxUJnXwwZbxeKqUOlL4F5pEIYu6sTjaRZwtJSULZVmhCII/Dd4ibSFvqGfR0wV16TzGHXlu
J9NFu2/TWAwkV8XsjUvp9RszqRpO3qTle34lCxBCMvpVUAhie1B7kV1pSQBmKPQmItQFh2jP1iAw
L1lf4Moo4097DN7Yodbb0ml3ZsZkRi0iJmuTg/srlgJ27IakTrKDRjoX80jGTJ2TVpjMAbOpWd/w
lEJBf1T69kZRpPdVBIqCuTizMIfs4Gnnc71cZX6kqKZJs/AOpYL8Y94FFX8WVNH4DBV6aKShvX73
k8QQR16ERVd/Ssx5wNfnPOMxnZVEF0WiixXYjPOTAhLzqPeLSxKfH4959cu8fpsA/5B3lmHYnczY
NUL906MAcwUVHiFnpfPHTpWaAR3DftQ8zXB2LdY8zKUvgsrjFH9Wqoi8iFL0L05KfxqspF7WoHNm
siPocV2Bzts6f0vh4jS/3I31lBT2zS/O611YbFiP6aQWchklx5YHJ4t6Yy/MzO25BXZFCBpXWSkC
KnJ9ZqsQmiXKZ0zdCBdG31k3ndAIO0CykDmn27IMb8tKEIJBy3eVIODmnotvkHc1TNxpOburWKRL
4l12y6Q7u9FebGUEXBc0uBmzna6b83nSi3aUCLoafu/OFufxmke7zLYoJXatHGosAo4nseSSxjn5
6CGXUoMG3ylQn62BMV6dCZCD2+jmE9d4wepaXYODlOiokfzaPPRruuV5LGr1mPdLanHiebMHGDuQ
MUQy8zp5lCrtFsj9Vw9WwjhdqHLc2Ka9j08ReDr8MG74dK6DVhjMNNjY6/dDxSR2P1BD0wnqChu6
wxQJar0odzo57z4M8fY4AFEnXY7fv8SkLegI5FDhlptFT3ap2AwdYNlFv8me29UHXu2wAqBKLxy7
IfyTTTz7D3/32vYzxtOZJhVegXIo/wxKiIQ0nRx14Ppq5IKb2Mnh/bzX2CKBcOhwQx526YgVxPiJ
RoAuL9ocGvutbGseMJZQ+OnDEhxNluqVhVRfDE4Ek4UPs/0BFrEtbuFyZFQoHiZL+xsDNoQhmHYv
9LnNAGSMQpzmE6HVvv9HCkFIuw0HqjTlx9sn5fQBQkwXrs5F5+oXGm10pHnUPO5FKcHJqliSsL/G
xsBcLm7qyf+NTTElnSp1YARZFjvpQcV6XC8B0Z/13qN5ne3ll4h77jAsYbb10wA+Qp4XY7nuV6th
YkHyZbcSwYcSQpy+9RFdypsv92EFBoOuFx48YSRAFVNn3jnT64iQzHgveEQL9Ut2jjZfeEv+IdJI
yOV2F02yl0lhQJNe1JYMrZxHVwehT9/KDvmaXlg15Gyqk/StibirWZxXbH4hvIZPDGV64zxjXHHY
jBXT5Q5UlZHqSKQFdTBFLdf/fVo23cgWGSppSNS2tCJLrkShq6OvWW+y/5mhicjv0vSRm2CNCuW3
Gp9VdU9TZjNcNjbXSeXRed7Q5iJk85fuwMBdfZODpgvxBbUua2EzJ+E8p8OXnBdAa7rYIRWsXIp8
ziunpKjOYxqMMGZ+HfgUGU6aY4TP1K1+FED8805WZnPFzxxbVYtzpzM25XBUf2W6AgTp3+sGqkBR
CIo0CkFsOkwTSh6XsDyneVZDLr61LO6TKT/SrYn3xyb5iAhyuW1mjln5Xjv0iQl5YRS2w+qazF2J
pAElHOJQ5sz2sJgudf9mjeWZxxzZSoQHWbOxTW13tW70AT1KA1vbhZXCZ/a7W5FuMJYXrzelYBkG
d2qMNWKMm+T4DPwSL73Kv4phzACbeUvrUsck2Y/S9jSbkLTfx79zDcT3/FTLYCcaH+2IIMrX+BfM
QKBXyLa6q+52Xek92dOMQ23VoQQgmoJCB1rcrL2MMoeLb/zwtlP3W911ELGQGKmCvuz59gT1YBkj
EzIJuQXWxQE4343TaT3sCVrtech8VglxkSPUuxwo4axUT6HrcRacKrIYsh1oBs35bo2zzze4+8kT
3iOgT8dxT9hn5F77w5M+7f/qlVoY6RmWgatDsccmLKlHQr0nHbkKvvN4g606CcuLME5FkoIb0KCv
HRPdb8Lk/qZbSbNDrNfRZOnKnjijwc5A0F72vE6Uf9xKyXkHKPudGcO8+o1gv3/B+X41y/unj3iC
6YMSlMosJv+NyMnYseTrrAmmz59Q6Qo8f3ULeg7fvr67h2QbYj33T0OPSqlcsDU2/xuV8H1v154U
61lQPAMLaI+5heqs371R116w16Q0qk/07UZ5EygnzRn2qxXVpcRDqIpiHbX+NarQU7qvC7p6cGRZ
7PrfLz4M8ZCtODrNDn9IzrOsYAOAd59f9OVTv5kit1Fu6HPHc1RLNXtxrp8BSCNUl7uumMVArT11
dcosCfcY6Ehz6nffrEK6dawN9g0Wt7U8Kdj6HzBA4OZ86LUMsPest7q6dnDhZUuNnAGrifbVFXH/
2Lp1ari0/hghFqlv5EX4LqONB7kMCBGE4zMDUWc2EYYsbbtamRxX0ADuKyf5RtWfyiP8Gm5RGw/N
hau1SBSKy+9jGi6RAAqaG3EVvSNsAXKvp1E7W7tmgQ+iRnyCVs/hCqFd0dYlXFmWonejf+/1zEs3
LTl+O7aLtfXd/XjwjdcN6ZJL47QRtjHGbbybUbOwzLQVkDG2du5J4QPoBrQ2suIj9MrqMB1Cb4vH
dFxzA+sjRRDKIn8JLIfVTcqkdRuXWurZ06g/69D8d3oTG7YGU/sSg9e1P/ahpDGY4VThcr1ovFt/
v9eXbAc/IcVyg3NWEbkBt+TVSgWRXoWUGOqC3IxCJPd1qrAe4bkVcAMIwbT4pNJ13bW6R/xCaBZC
s6fcACLrHAaiMN/1OeBhn/Zw56e0EhleZ/8lFn6w4+15f81p7XI5swEZj7BEW0zitHb3iJJ1UEm6
bU3ILK62+LbaQ8ZG55hfqjgbXa1XFaBRnAySQQwujbRUdoXiq3pErmIcW60iUb1pYDg4llE7rIpg
tMRcQGTJjW4RMetkf+o66sgSV6SysAUnAtFyRMTPkuI/z/P6Sg5HCiPyXfEeoHJnXhUcmqn4CkYc
Pw4/WSjH4qB+CNBXTrgFkSYxn8CgMwT+wlmoso762NpCfuMMhCtRF162mDQcfGOmpAa+ZvHZodtR
Sexg5gFobaYfqQ4lzxH+RWuWJ/J29lVHlnIjTx5eFCF8RLLiir3UzgLLdh1qbvvz7IRjqI8ZvjYF
w+49GK0V2Jp6i+76gZ1+EiF1NeD6zBFFermXfDK3seGfxErWCYHc769TwMGw54Nr/PPHxjSIP7nB
VFby8dTKxWdP1e7IGBnCNQbkmWWceNOakX9mhdZ8xrHAWhejkz1ocu82DoKqqXVsshQTA50lLdEO
QdoOaw8oGRZJVgmeRbCRV2Nh6tn+pfhyhULiA4BIdsAi9S1Exw28cdXXYBbZjEOuvpbhk9TiX3jb
z6TdHK4fXhRGqmbOB0W1uLxzd7Tk0ixH/vld3sCsMXxMUZYc11Hi5yimre/m7d12LJmfh4QtnBix
wS6rI175C8Nxq+zer2KpA4cTqExpiEq7bBywzaMbQ4ls72M8x75iWCnzG8GfGhd0cruQY+E+9CU1
V438ROJtx/FlUS43QQdUvdfg++XZNKgWcpjyr54oUzarUracfd3oC292iNr6WUbsI2JeTwisJN4S
vnzE2SRxMTVVlPUY9AZeDDq0VOD2ePpqvFrU3FGVhc6ek2tpcYdB0Z8/mX+M9tu9GSJ6Ej6BxsLi
3/ZGPmOkHC70LEjqpYfu5HRLDz399bRKan64GgtgHtyVP4ZhQVF3oWVXPHsrpRubaaXlFei3V/2B
3REA6QEEN7x7CDjv6yUpXwiKLkR0R4MBZiNHbVjXmxCJtTfn2LeCr5nfkTR0jliGuMQv/Y3++/8G
2B0P2vKuBEh9C8Gxu2KQHIXfGVjqZqQwgG5M4gAIFCaMl3jD5LiMvW60mPAUj56dXymQkcD+oP/J
ozJpmjVHp89JWAm+JTrXGjno9ChzrBsKTVfAZKK8e0FFrG69CNq7c0zs6r8T2somLWplvVneO+Rs
YlAO5jzMcB/KmPy1lhWIDA+VtBGyZlG9m3CAWnwBPqz3pNvDPCZChGXcigYktjq817CsGyNF6D4Z
5XGyfGIWkug8y8e7m8cK900zZGO/oAWLZJwXKac0LUZ0jvn5mk3DPaAzRw7mHZ/OKVC0etufLRt9
PE2cr2R1QbIWoMEi6GZ3wU3Crj3nzfQcbWqg6NHkTeyo5jortQ1KGWeIBMWGTNq8yigSpzmSuTDq
Sg9j7wktveafqgORhVAgZR4I6G1GBGcI0W0R+JXRTNxf3XRXxs6a+fcBU2s8JMRa/b1KPxYRE97u
CuMP1I89dC0vsaiymYgMfTc+ZOHmPnyxJRrG6kEjFv0k0/h/hSwwJ2dT9RDQZ6nrpzn7BHcG7FrM
2xQ1xSS1j5P9Z/hfrqVQppsRXaP2n+pjc6/+TBgH/qfSX0HazXnR8sbm2XlOSRNYA6wdy+NRgj9F
qRnukPk50bXQ4Y3tNyx49cIjn4pUblGwb2LTkMWhH4lTZ5rQSpu8KIFnwnaNUa5JdG3YLWZA2Jv/
CKP3nJ164juptfZW+h9eL9qEdL6NxlU6+RM+sAUXGZ82vFCeEp5wOEs4VPhOYLsrQuGEZ1gQXYhj
jNd9OqBOfREX7axbY0iheexoQ80xEbp81sB+R+Vd+Dvqs6XQpuLYffDicvRY5cWM0o6DkQf5VIla
ViMepshU8dS2zTno64XRal0UsJ8wSO5vSmVpYrne8FRA8Wm8bDwBI2JMUw9hSR2hY12/xVn5+8+2
49TsDlX6t38/0l7ofLMymXxi4pk4ccJjKdz95xu8O5t3ZHJnIGMq5Q3rvY173gFQra3x1fhAVe9o
XhTBZPo3NdS8mHAZd/p77RbLoq81mIudxZBOrbu9QnxBTPtzqnWa6A6xdru79TqsVo0q7ca6gAKX
0bCDzHriIiponH8GG8KiCq1pwrCSABc+VkLrqDSUcWexEDlRkkwBF+nli0XY+rkTYlxwoaY00bxS
r+6sSjdYEC8CnQF/Ymxw5Ci0Yn/hkFx/HV8Ppo9t2f6Y/47cw/vHRFnfsEVzhNB8aj9NNVwZQEsf
cgJuHjrIRTmX+cz2jPXorKtsIXru0atBOdBM+GeGl39++wD/N7mloj8DzJD8RLAY0hgRYLdUbbVm
IMsTg1FFwnihEn9MeHZDNL3iZCzRLCRCnYDlSfHbKB1qaOFkF5+diwyV9hRSGPu4UinXaGJvGGy3
uvViyQk+NX0HcRGWwVDt4/79LphNriwQY+l4KyMfP3wVrMpygeIpYDELJMtUwLLhXNUzLLruwy/X
vcQ0qAT1Nl8H1RaE0e3xceXYpUbkYfPwFS4/PE1FzT3T6/GRxh7znOJHKt3zm2qBunPg1zHpEXFR
gMhO+0dE+bCFnLYvjZMKlMIqJ/l1fVcoa2uL+jsGz3aELao2pQ1eqOqWGYzlitbAdlo3zc/saL1N
VGBSjfx9kEY6GskUd713Eyx2FM47V+k3QDK3JtBpAGs+RrOO/j6a7orDzJHnG02D7TDhgy49NaCf
ZdkAsg06RxGFc9hp5/QgrI8oe6ppu3SfbQYjpjvsKz4t7hdbNVUB5hu3cbdyTGw/g0xta2zKOOHa
tgULt1gIKazJ2w1nlVTtglP4UqXSTKA4VeDmF6JSX9+qTTdNho+ga01jOzJKzvyx/yn08UZCYnV2
sz6eKuB3wvP0Zx0Rl63R23NrZ4YicJtXHeYU5/u9Tcv0mioOj14Os6tCYpAIji1RMOTqUuXQufj1
kl+PJXs7jYNiqk5B0RXMC0phdANkGaxETmfh78qw2SBeFK8ZPJpDnYYb12qFO8wOkTjehJ82gyX0
L64i3PCkPQJs6IS3h5T0x31s0AA9KA5WrKxP5AjfPIx5gmV2CZsuCHHpmpnKvaOOL/4XvGSUQ3m3
hEOxC5nXCED/naYuppoWtLouPfBroXpX0AZFWZ5Z0MmLS5PvI+AXKhsYGEDVsZa0MKOdtQ0lNTUE
EZ20L/s7SZxQ7txz0ZBMUkV7HaHotZN+FRJYD8lxM3JeGX0hrw4kjubhE5+1sSuS/ILxmKBcL20E
Q+ENiD84+PcknymlACwxG99XC/7xElXgqhnaXBRxPf4tQY7I5KHTGS08mWMkXGpVDJFIPkyOdfqu
WN3EPB+0gtIMr6XuJ3WU1+gD3k9hNS+FkjoPhB0rWKrom4Vd5NQkxMGe1W0Y7fyx4Rpc/wKyaMBS
ryptaQZDCJpUrCzcIb7pD8w5RaPYQ3O05bhlgHmh8m0BQ4byy+vCN777uGQen39LPhu7OAs9ahRG
1q3G/IRwyooatf7Pk85EcCup43pdBG+WN9k8e1713Lyar3pDTkmjMatcH4edPPnJKeGmS9nXXAdU
DjlFF61zqIj8CPVpmFViuNr9bIBom2E+53gOp5Vsdyji2+8M9Zr5tKk93ABmnEtVqh0ilTOiXycJ
wxjaNlmLqqhogDuOF6OC3vi8zHriqSd9W90le4xI30Hk8EVsfXgocAU5M+igD5Z311wU5KWtLZ1C
9iGCnHqIWB4h7VW9qYLFDDLJnM/sqNSqi2XSJzJ3MeNGChmXFCuCRcQmyC2bzZiDca5GyffaDV+2
j+klm6kesSAneSt1hGym60W0+RTU+I6Z3S7L1LCL9kSVpyh6rztyVIWe3l+eNdkchUi5u8VlosTY
hiO4sDidM2xrEnsXkdjxEQsjdlCVwCcNbrONzrd45js3WpKcIqfkpPhUEVzPEwUOq5JdSaYFHwmv
h8Zu2nLSjmRFVrcetgZyUKr5McINQ/lrGNUl+Tnw2lzG6B6x+Em1SM3V5zgQxP06O1UefQNuaUHG
zf+0UHVp+KnODp2cnHCGCqibs14Ovt46nos2cFCyQvgsdX17Xz4tb0EZo3ZIVvRtJChk6V1S4o9O
8aaj4wMN1kTs3KH4gBL0rftf+9Dr3IysYYLs1i/zt/y+dHTnBnBqidtBu/F6pBYQFFRsJGT1af+8
Zt50yjmHegJnrGpze88mPEqYyy8ar6g0aNNQshTcMOlQM298x7mAyOzCCBfDdLYZRrJ+iBWYRffv
SxQ6D2k4UnpLBRlW+HkAakUENYYUkWSqUYgziI9aAICkTgCpf6wQdd9Hc6HV/hcloCITvnMalPbf
PcD3zXUbyeJXFUqM5pGpGRZYcWsXntYa08wBGqXaLyCHLdUFL3McYe/54lloJK0T0aC2/bxJ3wrn
pjk6YFdQOBcnIsTtseVC1FMYkfbpAw/6AwVUusyyLViTkifgDy7aXcbtKq0NXg1xJCmttg94jkua
W2Q7Ul+Xubo+39D8Pl0g9i+vEaG97E6+0uGqCveK1NrAN+S5kedzJ481rcyDv8NAM9IRAmvnHWPG
IUL8J5NzuifAWD770qrvO3nzUu7hYlgOxuCkNYGaGF/hVBu/ZhtW0MMVxoHL0MsUQif39k+hyt4p
avuYIh96JrTDNyZ0zAGPAgfhVJ+7RjWNXjf48zG8oTMenNuGRALYHxj8JQUctbjwDifZGKuBF9Cn
ZGmwFondgtfpKrUWXEvsx5soEi9lid0MklBJN6ZocUAmcuSomZwBfriAfggt5QxTwB9OlMF/Xe18
whtfm5LwURwxj02v/Ov3qNp3g+4o1OJAY1dankTQr+f4jCi4D+BNAis5w0TI1GoMrPIs0Q5SoVQI
zueNcE65wbKelge4iXDT8F9D3uJGi9o8uQ2EiXcqEv6QKJDkIvr1LIZQWaO5Q3KjN7sTYk21W+iO
URQXshltjbbgXf40Qzei+bVvxtf2ZmZrobFa5gMpmzQe73oKA9DHjZ/nKS22KpsyiHMo/igxp/z9
woyBmhB8oRhkIkm2xUGVLdUzQ2YmvYgJ6MD0LK0aGRetFZ7k5ADZOaG7DRzKhkCbiCgkunz4l0Ua
Bq9ye08zW17vUmukRGl5Afj9tRjnLI3/A9vs7YIlUljD55VpeZQeKwYT+rTAjF3tE99GSRGKCzmw
Jbr6yMlBrP0al2CFH8VZV/gHdJmUY8RDaf2FbU3dhQDzGf+VMwCDEpaqLWwpG3VVq7TGlxzg1Dgk
mRKX/J+W5BobzNF1QeYYZVuIaFmOMlvbRqDFdWSddoDD6xhbEwNVSxbXhZmc8aeqUnmKSitcsr7W
4kXLUGtYSwrt00ey8JteQxc+xlqsLz/F3TsgpzQD4XD+r9jCqZD492t2TqWCRmVWVxGFFe0BrGU8
pdWF1/vj/FTxEJotISzqVZgSRMysnMI4BXXmWPerKb2rTQG74PeYUhPIGOiBphOEMFK9aIQvry/d
7L19oayodu8jmdu9H9fwZk1Hg+W3jkuixMOZwfzdHWv3nxwfKfsu2dpUqjb4ycAyd+J+4fksPvZL
25ABB5q/Uct2KcHcz9zfXxllBHB74sSK7A6db8qb0EBgPxX8fQEGKML4oBBdGBX75xc64SXW05dq
n7RgG/zSsjyamf/v0aEw0bf+ya4s7A3o6Jv8stdqK5q2V3j32fejryZDPO0G2E6LJsLmUCHFrplo
0aSL5PBy9+JrI0SEfxz7Yb3PVKAe8pzouO4nNvmJo+f+ZWYvOQ+jX1Ixj91uIf8T3UqV8M94Liiw
t/qeM7keNDN0bzdIKkrd8tRXRqv5VmivYxVk4g1xLSjPJFgiovE6KAnPRx9+Gilv7IP6MvFbXe+3
v8NTv7ckr89xIsDZPpH7y1virAqJjBvPmvDP5dLAtnBrjSqkYiIMoM4UVgR6C9+UMv3CaC7JSCfs
3t4FBgZy/6Em7Mgm7UduHbJAb+LT30icszHd950gn39qI9KcIDIRYEKRqntt4ZzvyrkjygVygmKj
GlxTsXmDq5WWPdmzUu8Y3qQfgd1Y6RgNJ4cdKtc2Bqy9gm45BAbFhUdtdsFIrYcfK1RP5pY1M5yS
lQDJynYfwt3aX5v509Qm2pXpDS0sD07M3RpmrqC009wSIw088/VazvY6v47ULuQ8svwKLIALf4iU
zJCzNk4TcR8bHr/2Lx9UqPnAH37tWgmmdeJ61S8isKi0NUJrclmPZn1y1wCBUiBsUOq9t3m4/l6B
sIRfzsM+m2YtnN1QxzcrVLc0tilsmvEDThDO+OI/paz0tPihXd2nwJ3JzVvFI9gwPRqoemTcey0j
ubqq2zEbbD4PhAlQaE2MCz/4hjo5736atNDUNeuHFxHXD2R5HcCrTbpYGvLTXf1lvfDNz+PMIDVU
GYMXg4oWI9Wp/Ufe/xU/U+lE/IZCyLiApcZzoGirndwylQcvGOAe1nAp0spr2FMhI1kApJBmNBes
70ChoTH2qXdKbpbsDEHrbI44MZ09jgsNwYlUbZk7Zqp+/BQQ1xVGRwzVule6uM2U7kYF2WSCv/iA
qsOm89+sKSit44sk0WmSyb4fu2PIunla+fR/QK4Fj1h1WRfqkxzlES+AgtF7PMZiNy0j2aoKE1vX
bIKP7+8IhRdt8oFubgOsMiSRf3Niy75B+S6e9aMDApX3716PvA8KZ/Awhf+jC9JdB1DhG2Kxt8vt
YbI3jxg4EQCzZ+5LU5cmtTdhtklmDIx5bQtXxP+3+/eeoCQeQSF43t8u+IlfVLVF0aX0pyBw4INM
lqTZVdVvbi7yjrZEpQDb4X/wyU2LvwTmgocm/jLGl4/CDDUx2rYiHhzlkz7lUUyiUnRd/DOOcjxo
kqaeHZ7/stQYI2e4tgGnNKJtSc2vsfU3II671mNeZDv6UFEguA8eZl6FCnI2UkLK0qkAJpJuxBpV
q8p5rVSL7OnpIGIAV9ngZU42lt2rlv5z0QE22fiUa0FzG6k+zZWi9CRHoYJtgnhhrUT7DRLOQvJC
56MO8r/IU2PPcRCBvyiyIpyZeft5mue2Id+Nhr71OjOATSZ4/cvBR33su1jdxDExPGY5VM3EvEfu
kWf5Jy3GU3T54RMHYfr06ZwnzVyK4a7clDZu7bBcPhT+Hx3/QFIm9xlaK7h3alpDYevxHA+ZRSr5
0gN/LK6V2eU/sp4AdcI9Suo4/lIL7qOGNfNXhJVxZGoJ6ALXhA9/EUTcmQkV6o9vlDRxSDO7oOWm
3vwBmFga4fIc8l7Q3+n7Ln8hvDKVYtgmiN4GlZpwX9ASY2gzKgrYivFlHIKCITKTK38LNOI+Fb/O
rsAzqLXRMAANOZOx3MQmGIkZFpvhHVWOkvriVlWfUIy8+nI6F1pEYZQTYeI1n2hu56KqmkvuSPB6
xDiNXDSL6pDvKqTfj8KyNa92UoUfa0Y1n33vJnI8BYU0ImiptL2mdEokWLYAuGD/+VypBcVyNdUP
MHm8gqufZhP0l1+w7S2eNf3ZpJkhTtW97ZTtwlVOMI+A48ZzOTyJ0im80Oa+b05R16LRPrJpWkli
a0ymkLYb68Q8MBzPfQ51pAVmfSba1T09YINxK1rU7lD/ZuotsG1jx808mSmhQBKv+rdo4k3pRQ4v
7TVj6YpDYpCa98wAG+ZUcrP1i2xgjorC2awqukIEGsoLobtqJEvb7yENL5IdFuUhvRC95zIrEOq3
0xlBj5WKX4Vdgf9DljT8qLUjz1jnMR+tkQHu4lh9KLMforX/KEG9l2syx8yyLzf1vaU2GHzkD9fS
gB6MvtZ2OLe34cLGXRsAEKZadyHg4HcT6FQvngMzPb2F/fInxJehia3Fr1BrQX4p4HDB8FM6CkVQ
e3U7uDbXrRD1sWT78lv0cmN+wDX+pdMFdbtereD4vfe8Dypb6XuZuDxK8WxB7uLGzJAerWJElqXJ
lZBlb4S72299KHFE9MLAPByyx5U/cqzIGuqe7ADFD6JAS7GY4jyZJwGQORKFy0jDFDWoBaQe6Dv8
lBpoInRDxAB9DShdTmy1d/iyKqCa2cp4rOibjhUscXpOpQRYtMeYxDRugT/71GTCvg5EOi/C8KMv
TxJ8Tg45gNNWzReNoD+E2RP00iQBkzoeY9Zp1M49ugnPzrQ/uw6uNgJL2lx3G2Y+z2PTz5c/g41v
qWduDL0SfAwWwWSBtVsEMmWDXhL7drUnJKfZtee8DCcCaP8C56mbd0X96uB7mgSqdbsrIxBXv4HL
Z6P+C1E0rmvRj860bFignJGurL0u7riksWRciCvDwMckCs0SV6r6W8aT5Lkx+OrOtqVO3bkfxPX5
67wxAbHXBswG7TAfjwBrzr+gT8kn4K9wXbQYc9F7LQx6ECCKcEkYFiGDMMCxJrD45TF1yRBrJVRF
DrDfkvNsWSe/qdrfbu0b9SslomT9ra7vnzI09vy3lFfAFHSmRnIbxOK9ujRwbq560VHOuHDm7wsc
bO7+SAEFxRMI/edqZX672hS6S+qFSkYp/EoPCTnZyeVl6MUhDz6Ql4Acs5WQlLlT25SWIsDVLkmY
Yno+kWKzGcNC0iPaagni1Tec4QZbtGJ3JpKnXz/V75QiBxp0RgKBJ/5pTenxyHLFeuA1S0d2a5LL
bA8+Ya8ygSZYYD1nxG1gNjGaDQm6jhOOzRVaJMrYpZalaOU4FI5N5dG7Zmpt6R05eXfa6+iJP75k
jFRVKXfdRcNwVGyW6v2J4OZLDAbt5WDrip+PfhKldMrAxtdw4/bh9cpTNC6WUh1Qyq0o/boIASF9
IVjv2ZZNaGkErBa6DCcFepaB8plUz2aPGERU4OJ0An3bKqiGbsvAaWhraw2oUH2vQilyllNOUiLt
juMwckW5+2H2LMFvDDPEqsMQm/6SbqDrX/2iNwIX+Y0ozBv26omu+VfLKBcHY5gk9dVdZaxJgPII
bQyr88hoSHJO35TwAP8RCIyMkpDK27eX1rJZLoAM57dSdMFQn12LOTY58zK/h1AnZfsFXw44kIuF
1R+bsUvtUCdTGk4YNwxmDMOwBCdwVibWSFbWsBJHRazpl0myDKxSmikK/bHGZ0UnZnjz0r7bsSek
Ml9kt1Ao9VQVOP8O9Crz32Z9NuXOi9nqD8eafckCnFwJwREyV/cF4uwlftCcCzt13yjaUzm8Xto6
8ZMfoPbkN0U5OM7DTbhAImEcPaAGXL+hqKBJcX9kQeCMrCAD34M5I8nrszo/Fcd6fnsJoGLtVV6M
cQkUDfHoUuR8+rPq/hYR6pepaDeLxeXDHrY1cCUSQDeAIP5i9R0NW+IhPbdcEIWvf8Xo0B4/DrBu
KxAbE3UGDogPVzizMHWUHBp6CzhQP3wUvNxCRZcfDsBKxve+3u4QQiPUufcf6f6JjiiWC1bsii1T
rrnYOB6fsQcRabuhpgtOL000B9UAEWAe6BWYUXcVo3AbbKAMxpzH496zLk2BU2HSgCJqX/4x7E83
ugTycnSf2LASIUJNxXlW9kUhyRG9BbJrejImlNwYUVGzATE+pVv4t0haAa3IiqENYfy0/WAIWFcL
2wvWOnWCgt8Z6sR2RFGQA3Hi5tlkKQUuxhz6Y/rsSHh1LK4NxQ86OdnwWpqToY5RycISH0xKm0aJ
trvhN51Zngdag4eSGQKRYoU2Ad0pXSi0X/APNVgNHQRn+jjP8EjNSo7jaUbMQIjgvaBtxWNqr21V
3pyxkplVhubhLqF2flKfKcdL+1CbQyAcKA+eNI8JzubVcOzEMwy8a0cmHXAik6ezqgyQSSX9tN9K
2YqLhUlGnr5aMGX8TdYVTvJFLr2WpBHsTPB213G1CxSzGNgRXl629EdtoJwAoPUM72GQwmFfiYQp
tk7qp43H+AQYXeWYtpM18ksOV5/Mvp+J/VX/LVQ91UBNVqY8vPZWGIe2im1GIZbzGvNzxb+TbggO
X5nhGJv2bFviKbCAUj9PDsdrZQG1Y8vE6GIvoDNHncBDrPNAZSrtjVAB7wbRaRsBUV2GfVSvPh1T
z4L+0JCnImbP8CjrNIZqnWbNcamLYLd6yL7txn8hfJozv0QI+IuluGSxE9Sg+fCZ+jrOSrOsUfti
oLaSg80l/FJXHu+7A3CEKu6FhOLAt/O6OUBEEzBVwNiMLdDNawBlt1Pbciq95mwh60EEySc3S92k
sVMXFoOskNvN0yymBqCPMDxC3InPPR88syhE2k4C7AdYcDEKn3x++K7rKRBCMfUmXqithN5AHcFo
PpsArlVEGyThGssA6FasE1kJEHBRd5Ku/RYAMvIUDRfPPPZKSdYv0CSYPfb1NEbIQZcNd85cgjaX
JHuh+IMndsHbCAmUyPKtPcBk16IWltHkRZa5243jPi/nUX67KEWLZunCu9lJ2ffTunhpzXIugQu0
eiGYxTMj9D62CI5xNk7CB5mC+p4uU6lonW8NHHomr/M1fqWH33QbYS6J7ySzs5s9xhPj+F+ilVpF
+qdvWA/c33tPhib5OJfhpPwEwQLTHqHlT37qdpMGH3qkTploYWJ+JD1iZXyyM3lWRzIbns5wCOlg
eNuMOPVP27OTtpTp6eFqR4nCXL89yjhlQ1ipNdNPWtO6jY+taSJs4cKIUp25Y9MLnONKkqhgJLtu
/ucjWROREaQlJVmAMpsiPHDrn8ZzuJdAxM/RY6L9VvgkItpOHuReIF4B4hKyoxJvA9xIfCivjOu4
X81/1SlGBj3TtO6AC/G2eMOQ6alJMc3uGV9lnQ4W682xShTH6/7SlA3bOmjS+4uKYqk/LWxmkbVB
ydi9pRsRk0QNSp0jIDCgyjFPe6YLjde6cEk2SuosJwZg3DP7CWnyGiZknvbzeYgNXlhP5i96AFKj
IqBiBLjb85mMe69lfsi04/a5oM0tcuaEl6ihUHWxjpYYGUfLolWLXnOKbV1kbFndtKt6eW8NHjAj
jy9yzjF9iBgd0fMvkZYwBsyP2zEBBzDiSqyymz+Rc+igDahmSMglZ4lwec40Tt4cXAZgPBeaATHB
h1Gjtz7+06wdT0olII2eXQNpN9vGEMudZdA1JFUAeS4ol53CZIr2j3tBd4ekfnJtWVL+DCYzKcKB
YexcAelNwofoojbxPn2CoM2Uxxq3vCj0RfCem4wyh1uNpdnPmpN4tOoWzHPGers5xcUvvD9MziSq
4s8O2j/Rl/tpjQJ5qsV1y4Rp+/TOrEx49uCxSQeISX+vh3eHZLX9FV7YIyqjdfurzug1uOAc1yaA
4hy6lpECkFkvgdkv+HdK/wGmqVWIBkcZpxRL2Stf5QFY9To47t1+9vWbqegnpKCHzTAvg+4HobCf
XZaQ+AqVLsiZkrbl+CwUYiRdYzI+i0VBme9h40t+M8vC07AjSrNbCPGwEmQsYq8EoMZeng/nIPiJ
sC2ZggEvqMeev0SUH/aqhqdQjrv2HqH7PweIJZSesRqalcwJeEVnWl7QMXcqoZPnf91SGi4Q8EGR
/lpMxb4UwUuBuoC2LQp2YKyuEX6gCwA2bB1jhUjwJE/9kKBJSa62Ey1iaPk8qBZZTDLHw+TmnajV
HmYdaMxmOa7czFOXBZj+8XL7rQ/qgs0rAats3fiyIeZ4DF4ZimzpQevo1Wa+tiEhrN5QchgwrlZ8
AeGBy40uUTnISzgTsJBxHkT6O65aw1ypeQIYQlaHmujuNXcdUXMeeASwIJXhzMhk24Bp5meJHyAF
+ugma33BcFym2HNqoV6Rj6rCjemwArtUZp6ZJJSNPZJSn38I11eEb7KlTseq6Wsa/wCoIWxOmVzF
lNT00ww/domJemuY4KOWReQMI3WYVDugHWbkh/KNgu5dYeR+BN92SAynb2vRD6peE1yNeJGBOile
Kvd0igKG6SmztwBuQ+pubhoRhyGCBxuRN7TEZN5yexDE+ENhlm7JmI/oc+xFeGPiBSHSG6XiXeWO
/7jIXmCoQ89jcMpK5dbeqeNBz5kjpy+ZPscZNc2BSYTYU/6v0U+OlVnWu6WHtw+swvzHXxk96Pfw
YAWqTzQ9aVGvRHx9S3ZNHa+01Uid/UZMGt6mP6nqGUVWG3e25vFQ73V+kTZzfsSsKe9FDNaPZnsC
xt+AhT/JVUujKSh4y1jYF+Oe27GwEL8bu88reoJf2w3t2C7bChqESD9XuMj3S1+Rct45NAkKqknt
Z+XObmj4FDdnD3B7QkR6iQPBBTZFSRmZp+3+MBB7KJnH86YRowMffRhcjHw7WDGj5rqSgLiKRxRE
HACxmZ5DSVazOg69J0lrsFwhEUyACuMQk1nnihzVG+Xgh4h6snUK25K2VUsceHNAptJntelRQe8H
bwpR2m1VOIfLA7wAQqtk+Dw0zr28JUuaPVSwUR1/41EKkvHGmYbTh0FXP4JvS5tcKDWJkYNK44kI
8k73TxDh6R623yVIuZmyEQ+oExU+rEq66H4ti2Q3p3E2oGAsDKd2IYV3V46gIYmBn0MhFFTKyFte
8HKjOXnBt8MO2fUp2Sq0wz6Mkbi9+TKoE+ep7B4tR4BCLuPmjzA1O1hijzBUA3mHA6Pf1TWZnaEO
j1nbpZwK4M3r+f3oPZSxENpqr0CsXappoIivxtJDmSVgWWfW6cIN4LCfJRwZ3DAHK0cFtLsIXWMD
lbL4MSIu968JRf9OAEHzU+u5xNQOuTzRuFgnqqjVNEH6svEVk3hx0Uc8JEgehWEPw1+Sn1de+6kZ
2A72PQ1FBbsyoHa0FYKB1iP4g2zigVerId16WEyjUfxuGmSuMZM+axv6z5P1hOFCOEgzFNbzuedI
Dg2aHq0IA0nm0W1chtmD0wX5dPrY1HEztf+LkJF/vYhoM6im3oQypD9cQspxa+tZ1D9anf3CsqN4
XZlLhQDJEd4iObGJ/qpfUuq/zlm1LzYeC41kMSoodw23pCLMvFcGToI+bJO9oR2HTYU6f2+nA6wv
Q4dsowV4+lUnUIYMnS8mxRb586te7BKwLI7o6kbGXRWE26JKVWqx9moXfN6BsAr3pZPMg/UaI+jG
GROUEuEI1/54MzcdtB7SEaJeGxJp/qfd/9EJMjcEQBmHIz2cjXG3iLru4ObTJFUaVB1Y915t0r2D
UweW5jE08dBAjbxfmv+eiIBZ6EbFH6K02LkeLlvJD+9henthwwWUBJGyJ+/KGaGzWlkiSx0ybYkt
JETpNeSXZJADS7KMMCXbwMqelhPFSbuWjjrIDHkQAui2idN2km3TKaOppRI23Xq45Uilw+tj6ngt
+RwmG3UGxXHoiNqKjHIUuyfV9ljzK0PXtehj8aMU4GJylL5jyYB5fVXcMvHNP+QG7l/bjuHlsNbj
TELz9VTQpX/+Xh1cc6kfsj4kc+KOP3S2FDUW9B1mSTFmv0yLfdgLd6yQfjGT+cm+ETBkym10bp7L
w0IcyWiwLjuQHGC0IpoF7uxk0ixrteRxfwBa4TbPbdNRnVOAroX3683lkNvkfAW+gm6mb7KAYirR
3zpugXqSJ1E5EOSUny37b1o+JCEVqAJ/y9joB7XajqTadLBhFJVzGk8ABNEH4leYrl/H6c4mYTqN
VQAM7kjY53SF2SJS2YoIQcCakmGDUpcOjnAHzQifS7CuKOQBuhk0c0IwPfEy+4kHeLB0PlmaQ4up
kDXlLRTRZKY3dZeniBOrvDTtjEFm1qwy9byCNLdleoE2QNL9mDILI5WfIKUlRrnHrO/r7FzkdmRr
cFb5r4HGxW/K4rkZuzolKvXMW5iO29PKK1zGfGp4IKdBfOPpZz+oclVuhP/tgF2V1nKHLTi4d+Z3
l/eF8qovZJXv6ZjpdZrbiPmM4fRc4TjwXbJEFEo3FUdJwv2l1ygXi7TEpn5LmTD/hFUxZ5l4e65x
z8d/BuCFmxk4tWFwejYQtxdil4ssBpMkfVkfVhCeB04crqGSC/i9hcA5lAQgn5udg0lDVlCV2/vQ
7+E/VUE+LkGB33l4JKsMlaxNF39dvF2/pWj1JXBv0Nldcy1RGlrl5PSDoGdaZV73GABiVIlFs7Xy
s16CjfaWNoISoqM64/fO7x+5y1xk/qqr5wtMHhNF+M7no3LwLuoE622BU5snvsYu1wQPKPVifMPM
fuJgBZJFwPwJXtUb8R67DiWWwzIG0eDfrtcfpVguuxJ9uMJ324pX8oN3rmHe02rs0zLnVfvv+Xlw
d6hKuoxNGCOJqEqXxTdj15rIYXft3b2EWAKzQ0a1Qo4K1mogqZKCHtb4FCC9Ee8sB1FaKF9LKVD8
iRDwrJ5YWRGafq8iXKA3OlGEvZFpG0UpVFoA3KEqlC+a5dDMozecFMRfiaUhbuR8nrwcpyqwiUUB
YH4IUamRh+w3tKICASRwPtFddeqSGznYycZJv7hDXCwEsxRcXxQrY/cI10W4Kx3zAfCIURKtOEAk
lxJy7hzGZHhyCmkt4MZq1AXdoH6RS4RjF2RR+TFUbt+IPXKPimnw5k/SKp+NKgG6PDEMUVFLnEmn
WhPdzyu8r+9ar5Oa6lyYUhfNeheE0odxn9UROLVweERAJvvDEzFGuDToD1No9G76U7YQvuxWT6Xz
Z1uHAfoI7eshtf0SgyMh2OP+Ut9ZyL1i/kRz+JcduixWX/+8eFO999GrSAwbNKsRjAoUkrLxb7Ab
y08O0uRJgSs9XEXsmSsts9tit735e9iEIdirtQAp0+2oHXXlgkCcJ1l/niCJvg0UbysNIvfhYo1J
IDKvjDXmv++iBl39Tfn6jOmy/aM16iwUgQpUMHEVfNfvLhBpilsIygWRZN5L75/kYMtUJCjC+J0K
GDmMv9EC2vh6XxfVwVViTL62HahHAms79TOrks/fr01V4L9JVRUyMIZYzGLSZ/pVAjTI5c+SuPVt
cvnXrZyiqbA3oK3eTt3rPO+UjCzNjZZPfKme+FeWuCsCnde7UL2N8ZmkNQMkPhpL6bD0eGSaymUL
f5BVMoPkarlxsqF/Y4fouZ7LeGr4oQkQ79TS4QJ6UXFmR8W5ox3SGhWloz6Pj/Oa8ZaNcNe/0+tY
yN5KG/k4CY9tvs6yDsjNF0TJvr7K15HWZawypBy9f4Gc9bGYQ74YvaacLtb52LhozgVcwebw+xVy
DoKbnDYYyv7WNO8ONAazXP0xC47uogzxTVP0MhbkdA91XMyKdiTADW1Idp9YQxdHuz1bOtzNCbds
DvwwMHbzupi5wfosHVZlz9emJDtHbztXVulVL2nh/w6Em0p3ALhs48f9JesPZB49H7BMrHtX6dT6
g638+wB/PL3lFuy8bwMIbTAedBAf1QfUwx01TyiTm31JuEiY5RFeN8C657X2xv/jD29+Ur1Df2UB
ZQip4MBuoH4Z26HNfQX7uMJ7dOq5t8txRIKG73E4x2mHwoLDYZLDtsTVLfBSnU0k+0Cv7f18HwcY
29lXtSdLg7a3cLgmx+j6fFxVWmkYEM39VIRwc+qQD1ZGC4PBcBqiy9lN9QMYWqM53fFtP4iLg6Eu
gK/at8hoicQsEXKQDajhrHg1SkviB0v0EwvObjUHPee1+kLKZNbzO+JhJO1Sx3lJGNN/nrzlUL/C
76hieMuJwciK+HMvAu4+y3X5nDBR3p1vbqi+nWDor02kPCYhFhM8pHRDWT/3ryeRjc8cvd7WMeEN
+nlM5RiyoG1jHiXl4TVkIcY5m3LIcv77T9S/O3/MUKEqrgn/i9c+IvAWE6E2Y82WGjAPVV3ibWGd
7sWXGIz4mCwJLhScDW2EucgbEBYdAb6A3KSNvmFZT6aFX9C/cPfk4TfIWQXd2+Yxi/93A0u9sdAn
aq4nXQjAoeDuYj5aB6/69N/jXvuwZc3tjI/5NGTs9AjQ3g/ChJUScln+IEbKqfumL9b6JGDP28U4
UHaxj7IPc+3yBcKHxqGBkDQI+8zkh3PVAZB4fNdCKN69uZIfNK2UhRkVrimder3CM3+Xj4wd0zxJ
A25BBpp/2Br1L3mmn35lGcimMec4YoQ3Fk8DEU1q58NTupmvHhL4yamQq2ZojUFVkzKCF0msXwEs
EpI+Earn6XnTIzKHy4ttrofyPGbkKiolBa6DOPn82Qhu3/Hg0TzGhNXVfRMkM2h8lyScFZ0w+OdK
AyMDjYdZdcpNdRSUreAuDB0c5iKDVKN0ILAHXEiVjt8frwseqpbbjvaqbrpWXqA6bvDdSRVNAYvF
mQcpdewiwB8r6KxugJYODglK+9uDaqc0TNa/49Sy3tbzefWiPZwgTSUU3Zi9JTkccPUoCcphYgUt
K0nYosWUipPi146ugtDyxcsz16p24SfiRYPhEhSjix2AygwHuOi+N1SZVde9QyFD0SMspMVy6O2B
XwnmCWso9K3QZ6+4KOFEETrbGsIf9zbnz1rNiWtLYLNhRloTKBf0ymS/Y9LxsZDB6wm7Iit+lxHH
MRW/rXu82uUzue3AmBbvyRHScqS6Gx5TeWILZu/nl9bHM+oWvw59BcXuy2DKO5iGzkyfAmclQjRY
kqn2YqQHPuig40EbwZ21xPffP0aeH7/bA1oYmwC8GDL4U9D27IdZSWWPqDZ/Zh1k+Q609aqXeAm6
Z6F39cdbC9najQ2gQ9cKsRLkWsGkvwEkRcoHE/Q/H4seJgJsl48+SFtoQXbW8t4wouMHmccs/oBD
dXac5wV6bbD0KBpCJknP1zWJB/dVT8ynR0jsgQtbfN9Q8d1uVuOHX9DkJhowZzpHUHXVumTixyAs
Vk23rFqcm0QV1lX5mJHtwx9JXGZeQmzAgTj37epyfOyylLiWIieNU/0NTTuOqCocHJhfYkDbE12i
BaSfNw3QASKMQIHgJH7F3lKp7Oj9rILva2hDcvQh6gV3kTsmWKS/kteJZhoPK3eXn8Ro0Zey+nDI
FzjYwRNE2jB7VwVpOR0BSmNoUBOg7xGFVgtTBnIWYjOav/6GnjeU+gLnYfTeSlVSLAqgncyYcRzg
XtdmRaRpEEI4HzoEzQBZdE++2nsQfhZcqWVgSCeiNCh+jjDAj8pH6yHIAMf9M88ThYQPRNUYZFxz
joGokeJyBFa/ATjp+3a03B9rLkECz5r0noxHaUfzoynMVLZ8Lcro3RbGQVTIThzA/EC9KxsrShHl
nZNFlmdsqkEjGlz8yV25fDxXsvexL2HLFRhwUUQzN3dn2KTY/7rKpvImUHt2k9HyRNmGAlPcIJoo
ieAn9RgcI7uvapfSE+l8AIyxZwMbgZ0A/mgLtcbwpWLUN7+Cek8SFjw2lQVA4Xr1afTwLkZPsE3s
pSKE4BaYDeAPgSe4LeBQV17x/F8JdGX9+DRqi/RHywR3oTlln38gRjcY9C0cXsszEkcDmp+ObnW5
4JyBfFLr1PJVdHN9hJTj5TH7vxeXNp2cr4KOdDyJYuYNc/lVvAlzLuNpPD5Miks3XTgoASd8bDZf
NNc32dIMtzwMzFqQDUS85ELx7hiuk0cUpLxT+SS5YmQsF5Y38cc32IMRHMcAfSb3fLKbmcrm/Kbb
aL/+9pMfbn6ZgNq75kEpZ0Py3HAN0A3cEYhHvVOTqmKqW7jvMi/rm7lt2Dk/shZMemgr5hLfIabH
cKxAPP58zL+iCTrkBWDo++PVgfaOnl0owPpSnegiAAHpAGkbrJo5HXfnf5d2Sy+L8s+g+PdQ9Y2z
kvWmgZlJd27F29acPjZqzk5dpf78ENcW4qoZupLpvwKTUu5v95Mo1a3xToCsWg9NbEkoSBDlyz77
qrH257KUX4XVY1SLmH0h0q2WHkpNxOtxJME2DJoBjyUlCEPd5eDp36B8I8nD+Z29OzXKpnDlAtJa
p1V3A7inRFLvZHqOmBYSYRVhRaeoGgVZMkaIBNfRaQ1CBUWHa7cuidkTvkBmUm2ifgy8QQh93I9a
ldnkVBiOS2F15ih9dacXL1uLoqrixQe4j/gUfYCblQ59SniujcDE0/5popq3Oc6MMxKeKdZIIF8L
e5sLzHWcF46oJwhAPElH6aCZi9k4NVvykn8hELn/cTJyoiDLZhg4wZQs9onwaand7sUzCVz2aKo0
ypF3bKKBzPhGygYZ9gSgbyxKzCQ76OeL/phbqmrZZbMIeVWZ0yVNfKSqTT0iS1ep85MsEFO7KQrU
OhZfsba3wNOvWNXdTswQXwQRTCcrPlTVVwuN97lhJIkbk6wKmB5zWUH25lxjUoH+eywIGTIbNb59
FhWqynlNEElHopbMXTv0D4dxKwtiiYo0THvi78oLdBjxu1bewVMVjuXERpYaHcf595lTbMWNaeLV
lmVKufvmPhr63E8n462+kSPDKy01LVuTkvR9tWjsFbI6ZAAHoN+CGuibLn7+Ik1WAYjNF8S53Dbb
hg9fDl7wX84M+ub78t5OBnMU0f6bNKXy5O7Aep/1I5+8CKhZh1b+/pO5vExCmZXuu/PoQ6tiZnwS
Mt0pVcPvVBpuwDOBzdDGe4mhlp7p0tgIDJSkQV7FGvjkEr5PqMlKPr/PpTuTkyrisZ9fvV89IAPn
cTmbzY8Q5jAFXWV8lMDU/qcTDOKI8nAmxZzEYIBM9tE3B2b8MdbxZhDuLJICOQQBiKKui2EhC5Vo
haY8dFNyH+AybemQH5yZVDPhgvIhLxPRyCDVER1J/79dvN6PLJmikvH1fJJ72UqOe8D3XSQYPve9
mwqQyq/1OHzAX0YfcI7ON4M2AVItiUKIwZTf3Ygn2mQF2XHTcS1UgUM22xjfmBk7ajQSN32pwOIn
w19JuWxEA3m7cQZTXCC1+4NFZZvYhp1mDWdScyWZQZUhL++HcDzU3NiKob1/n2jj0raEBUeCLHFM
72cFM1UCDoEsVLcrVtABwJx9KT7IHw6O1y2nDMEkTQJzcy4qJrlQJPsl9nof80r/k96dUOrdxNQd
yLZrNzHwF3HcQgxnr5V2ITpu1QM2bcGForwqgDIzWTmv/Dvace9iy9lB1DX3dFN96yQSMlQbX5bC
BhRphC1LJoXHzLbeZ/3tkCfR23hPJcFRXzeoTV3qs3yaUEsTztBryppRmzvbsLG5FDt5rAk/fmOY
Rz0iHvKQX2DGUsrOtuDkob+l0sRZVcMCeIjUn/SgkV3H7lRn0tDTBjDMOgC8t/9/zL3s0jCaU0Dh
jLrokWDdBWEdtYvC+Q1IXZ+pW/4QrtYeasL7LQuFKimGe+2R4wl/6w1DIwLHchaS1qISOhtgBFIM
+1RdgO4SBbns1BfKzrtLctWzpwL+VXGOdSnmfwrV2h1cPRXDtai48AXdkpOGLyCYvm+ObW1wh1eR
TVMPeqNEJsvjyLePqC+Bbv2RH3YHb7E0bvnHcWxO7D3BrmZFgoN+TR1bgHhfv+qHIZxW/qOITFMz
B9u2kANrTf/ly3t6wlXgIdLm7eJajju7VnoWsqjM43dhSBvWrG+GTDEyWjA/+UudGS1eTxPhBGD1
0QrRUOH8oZNqTs2b1mBb6OM3IBSD7Y2NnKa/4a+tanefTcf9dNpQEeZO9OUJpxuHGF8EZ/DoquBH
bRizTc3DlVQh9AIpuzqxQjosGO5hU7kApUVsgJu52IU8nHEl0KylXk0aDEs4IoarQXVFEKa1C0rU
h8SB1CywYoouBD4v5lZzUUXnyu1YvSH75pQiFbvGvXHVIWT7ZT3CPLjYKtXlXWnzA2+62gxmEENS
hGBDYRb2lggPfdBqWM7X1WQImSmwQSdhuAiXmRyeb/NCxQp7/LEyqfUiUD8jITYwXuGtqsGaGlsK
mCEv4oSlHcX+68KuVOyXXL4ZzhMRRMEXyWNPIdvY5MQEvsg240FhT2zjAD4htpJ4vFd6ZKlgRfPV
ge2YPiF3Z8QZB+O025vHutQMw9IYtsViQNQ0X/LFrxJRF8wd7NVaBWpCu/TPgaWF4zzj/F6e4qjQ
aegAoVCKI1FQBrQanDpID4VZtFcQleh88VQ0CleraaXSSXWQdrWLj/TF/JfosppWTNdXnvJmRsAm
OdYouE69oZUeZx4xVNYfSx1H9BPwLtJfyOvXsN8K9ST2aXLtr8oa2bLhgkyvB1LOrpKiaUPZOFQl
mW2+/T4TgJQRWeOZN+OM43Ox2aPspq8GxdKPtOVzZY7J2IGM87FTxKzGJL0lDeWRwG3rIv7Yolqk
3w2g3HQwZurNROBqOxST3PynGIKdsjAKG8hlX0gSOydXDEVUjtUq21i1TYh5RBqSZEptsP0vUPDn
L8QkTNE7/bFdSztR+r0XsgReb/VdQZUD2QpkxDFtr+IWUSLFhUrVsceukz6VqZ5BvQZz+m4GUEau
FXaDF4QOfb7biQCkj3/5c4/KFnmyVGHwM4cjVOs5cje8W+X2vgHJYlzhj4inC5TU584CdsmBBvV3
lA91WatHwT4o6apyuxugArPamlSNsHO+WgY7dVK6d9HA6qDqbPlZ6awOwyswv/iIqpMsGJEQ9dqZ
R7kEUzv3qF3v1NA80Y2Em1nY7IgeR1hQMKwL/AQSpLSayRKC5WEQYjmdN0+A2QdBikLk7u83XDZN
puYuGtR74Wpn+k/tUB/dJwfbXuGxi+vYOt69opBVZq+3W2Ji67scG56WZ/xCF48yS6h/zSBVlCRX
yQnOxJLwMacJDVtl6zQuR4UHAkoPJgGezgthxGCUHG7OP7Lfp9MJfUXgQu3/q4ZFcggzWXGWvS2T
9TU4orMbgGdvHZOWJC5df0uW0dPQWxYXFINyFaetuKfZCdtvgAX9n4d8JseFcPCUcYdT6NYK7tbU
oPg/iAVGi9bxeBWWJOWOZ2n1DCW8sTERNQeiT2gSDv5ZJ+oMZeTxnt0m8+NCtbSYuWeSX8UI36SX
6eiIZVR+5AnqqZ03F7au3lATBvplRDDWLUKddxblsOqJw1v+stvAMaDrh+J2bY7vIaYFaFyfkJ8V
nSyfXNuSgliAoCKgUbShk5cLxLGaH1OKuZjSjJN91cPU9JBO7AHFTDPa9J/l3RFs0rr25L0Ax84i
j7WxN4La6RlhCc7BiM9iHHBZtbI8M6KC0VKUyq5m8gojS/EITNDC1b5JdG6Ub4qDnr64RuVczA5Q
mMTlZzO23J4L3vTlFpyXDTGCrVU6PvJAiSU5aYRKGWmlNVtXn/k/YEBXAbatSWnpH86fCML/PsSf
bv5NUn7Q05hxpp7kgM7hdmXCLvmKFpvHFmYIZETPFTXhxCbDD437yYYlXLXiTRom9qHsYxo1LxR6
NlGHd0SUbVHFvytAXS99uGfMRemgQHsXuwDSEal26Up46jkcT6firjXfnPPi3y4iguSpxo477u3z
+RufdF01nlq9f/23peTrJRcnwWCVHY283R8aDt++zJTlvaprJ6IFxEIHlCOLfWUakUb1LtjpVVvn
tPprNvPwaVrI1BVNKeUOjI51PFeIQ6X0bqJuJnR8mXfYM64LTL2Mxh9ME2XETKShZ73uR9m60D17
pe20xH288F7fMax+2M9CGHKn2lEyhzlMzWnBfOo+FhtdA2Ak9lNRdP5f+CUsKITInn+kdQXc5Mvs
3E/xR3Fy5OluVOSQkIXOQAuWurQP366js5x8rkQJG9jpreo3+zwFsM32LLivQ0DqrjbJfuWPsM/G
Uet/gmRsYwR4JDZdV7A9pRM4flRCjSDjjAZrsJbweSTU2tt75vYyoOvdHituJXDouU7ZJtivuFyQ
F3594nY00oPYf3t/piVBKMC2Xm5FRWnjgXjYfwju9U7PdpNbEp93ceyT7JfenJu6dIojKKPH8XH/
KjymglwCbfqtt2JnEcbPUzcDAhp8Y0AKnHdmER++/RPRSm8FOSnJokiExqgPGg7WbMPIjnoxlOx0
N6BmzMOiFP+V7VSVwpZgcdOL6MidxS21T6RVfVGI0+SXbqJVfo77btB+bEkMxyvEMT+CZQl2L5tf
Q8PKe2d4fjZcI7FmqXNVBQD3h0rVGgh/A5Qa2xDT2roy9B4w0kMtJ6R6z3vJH4C8xRbKPn+kqMLR
6bma6eZXCSFWUYS8FcSgFSD+zMxst0TYrX2SI+su/10fKz8Np7s/q0EQBWk7WE/+TIs0D3IODULX
H0SlxFgoERSDsJh/+Se5TrzfydArNq8XOzzp0EnZ2a+wAxRW+or78Ow3hyKXOq9i8msxLwt8zFQL
R4zjXiFS4vVJ4UQIhbAI6dDNYtGfo0+kQ6kDvCUnaMvJwI6gasrABymHJdSVHtRypvATsWOWtIdB
mTnyEyrWFL7MS+1O4ApgFTmDnbEDzQf16GuQiny6p+CZwvEL+9wxaUMy2POzHA5dWasUEreGOQwP
zfWKYA/f0SXRVdyl6XKtTe55vuegxoL5HZ6soIdm+YIGibYtBkBTQ1x5ANYsS3rm3R+Np69um9Xi
spyjLcM0pGgNzWLgbGdZACCr4aWe/jmmaHptAY+B7DTWXONXciz8G7mc6slUTYc3idRmP9q0mhTi
FlDd+Fo7xQ7F4/8UCOqN+AJNi8MCvn0U8gesjz/yO+kXcWYOg22MT81Rj/F8tkTeRj8T/7DJdBLw
FGgD7iJhuV5KbDorUppCPx2EBfgmlnCgPIMGOWzndTP+u6hqDE12UXBrWtN5ISd2i7+AydsJWTpt
q0dLlz4y81K5o3kGrLnGBdox6rVCuI3iaguupz0uRg5MMb54hfJRumvm9uu9e8jWQodqLBD9+Fqs
x2AJXt5MzdDvf129tlygr8xGz5l9WSFR5HN0wHZVUp+eK6lMpjhsx/U6ujcTVxouSw1i5pkMk98J
uuvXBOm9aBBcmsboJ9ilmmFwqnz0Dnh4m4crjFBefk+NEUYhiA47YuZS+I3YZyzuN1VbRx+WWS7y
ucv65/R2h4Dd8jXeGiYyn1Y/LoIwEyNTYZPHcORyTP++nztTk6BR1mkjsf56ISw0WxSmvR8ekl15
lK5r7JqF9KzzdBa+GsCIuEqXAf/CVWPiIeiMa0tfqp3zcI3XUcdZIq2Qd75JySR5IQSXIFZJuOZa
0CJWoW/ktZJSfyv4pLraMYhhjCdRiWeJgcehqiALumuG3BsNknWdQOW2Uw3xuW+0VhNK0R9NJxOI
MnViKNJNEyZOJ3UaFrpLQtHTrVVzCVruQgEz+qPVB0Hp7NK8+KnngtpgdmLvCfkSAO7N9ws1uB4y
zPAb9fGtrtdPxXXR5kKx1wwtjRTRkuAPzJYgXtf6u5bXjpviNnhmlDTCB1qY+ALq7YIcBx55YC7d
OnKCEKyqLR5oeSG/yjzLUFdq5Dic5Wzp3gJGXc/3E0efNPEueSHc8f2EYVfiG9rPGg188cTw4Mf+
WBt/jLMTTsKVCuKTYH6PKMY8zq7AlnENhAkhRsRxCr4gvyvinks600XOy4aoeafFE7F3Oht9y6Ph
mNa6TxPshdjMSJJfrJCjZpCuw6ruZhxwW4CXHEnxGJkQb5xzM4DkO/p5q36wlayg68tOjqg6QsTz
Ib4buMf3AOpVcS/ie/7Q4dl2QBg240Crc4f0cAOb/715jnTEuubMsAstidcNyOBcblaKibJneeoq
g2/8oTUfTUqSATg6kyN72NtvFcDuZJkwCWkj/wu/VpYMcqf/Ut6RuWZ5Yneb3VFyHQcdrScmgJ4O
z9TbeNzEktlNgarCuEVe1L1Pgwhpzbgf4EuslcNizSQSEfq93Qwulf8wqGcDLKVghA73U2YLDgXW
/Jqwc3smbMpi1q6bHO6qhkgK+8XnTGWvQ1Ib5qAnbblBSqacikR0yFAz4457TlIL/TRwdjWJo1kH
gcSz/Fo/AVJhhYjk4v6LCnJisTmSgG7lPTOaJ4KxSrPXLE+FYz3T/unWWEzQJW4lE+5fyju4eTw/
G+q9w0W2kkEZUc9riSw/fT78La4VoWn7p2jk9IbqtGrDadOBcouJilOR4AsSxKDicAVBsaHmjjrq
Cdr8QN0x0WdeAh6r0pa8MMHH3YzMFVaSY50tJP/uGJXI60Nv0TfHUnYvQMcXkvBOunACmB/JNt7l
YG2FkkjtIqepP51Z4bSJVGVkFpEqK4vN1xeIX37ZCmyJ54J5S33jhps0T98Rxp0H1gdyaPagT83p
AQGrCsF7ctwJoyKMUDfFSDXaTfe1zqe9IwUGoRyjMrLkfCx7pmn1Ydhh4oJlbyEQXaQtCH+WndjX
xHkoxybq3onsR08qY/oRsJQobBJMR83P/VRtrNi6tbHf/NzGq1zsr7fxxFim9MiDIV/eEkuvo+5g
bNQIfRvuHup6uREaBsws4uo6i3WYwFln4FLVqO326szV2yOVYnZDi9QpHO2RAJ6Yl2mvo4nyx5ge
CwmQjwKNMHCRJf0SWN/eY0Sg9hOel05DQlVdCdR3utAiyludq15ZNWMFHOJRG5V3NGNXdBpfAJQq
BPRerubhUxuQMuki26QicVggRNipB1tjCiCahup/+v1YqYnhXsZaR9w2VN5a4M5VVBLV/FE+UuQS
5RlzfJXDKDWrB21NQ6UYx1kVaE1DRdsiOIUNVMbcRpF7N9lrbZjbauKCz/oRGSxKxd5C5bdX4kpw
CDNA0xh740hp+n9joI6izO19e6m6ZVsILd1awzeBSutiR8o/SGFylXTFwutDr+BJC1GwGf0iCqih
yEMTVF8WgSFFy1/AhWsYaxQOgI4qe6qVU21NqH2SsLFb91aSxl6P3K3E+maAy4iISInAbcBu1y/9
YHyfJXsEz+jQlKbRNsLVS0VOxBDUQD05uAYhc8w0r3DKl/JIcDRTxtqrhbaUsrN00Va7ii8iHxV+
zkJuIyv6rXi4/4gA7CwFlfx2QYArRiGopCWOs76r9cr6xUG76YITE0FuO3XcfoFstw7N++YQeS77
fH1Na79nHeW9kYuF5GTupktRJ7VjXaPNjLLXuq9GQyaV3FmJiTIlWchvIX2Y7RsoN+x/fkRurNMY
g8QGzLNIAMgMabb4WghxG27i/NbsuBs4xJKScOE7CgCwXshO9B8nETTtWekZhbv4Gq6XAmqbsnyU
+vCj0sUe45zeWtQmWUS1qFl5xjT5355ofBP90+MXgib3v4hW728yJZaPjuXbEgukMYFRSNGWIvlF
zMgo26VayeNIIYjlf7kUKPzKbs5JIru58NxcwUaKrVzqjKIhDtDZf4Q+Bk8t7IyvjzjRiBsjEUh4
6nR5mIJzJ9C7WJ3nwerGaKVXtxVzAanV5AzEJJa/Xnr6XIefdxlanG/cPD6bTDvVh2eYmeNqLWsR
yIaZzYbR/5yMTliXDAPfh9AMAtS8g23cq0Z26Jg3PPQZql4rDbAwROuXrd3v7BIknRn56vKYJYXN
aML750TYiRcnzaT+LvOdI2VEQ556pvHOMdpWzU6YK9FZipRYuWg8rYm0WWJSAYF8Pmt2Jo3xT8Al
Uu8J93h7clSkSTTZB33JFn0ohLYXTh+MWXybJXLrcYM6N7ACJhqAE4iXR7zRr0SF7ZYgWYsTf6Je
izwQVQLCHcxvPprXwGS2nGCpRzy/meKDN9DDjJzw+SrDs2JeiICNP/QmqaBxcb8inxHCgV+N1LoJ
w9z0b0wJ0KFLJilbc3UeW3GSDlVWIHD7wAbf8vFL4WxfUlE4W8Q8BDnLsizHvA9t6WyCgI9E6A4m
CGOsHOvFGj5c0JIwYUyZh8Ja6FAqDm8UxpULgqg6K6lzc86AUCUdHBA0r09TUfuOEm3KmTdzE1vo
fsjzBU9W/6vUDY6SMUAQUL5MUqrgU+oJHiYdS08MivgFPqUN5W1vIipXKq9WisTm8zzVNBWkvMAX
0UjriQEeAbjoiCzoRB74ol7r9s3hANAtyxf49hACoONUN7huONCsxc9Igcw1kfDURWZjkXes3pUs
C4TCRSjroTkUqnbhv0sYWYzgrMgDbVxKK/lOilmQzn+rnLBhes5GxF3jpvtM7SnIZMFPtK5ZV4eJ
Pkzu0LZuzzT+frla8IilT46C2pnEomsIY69euFC/P78xHGBj2Rr9xqJ+mC7jTXoyoG0jK5NLoEH3
saQ7RN7Scc0U06pr4WPJVOtmuGnVeisKD1z+aGMjPYl4TzEisORpVJTUt64aa0iZOv3m8PfZeBHt
avZxL4Crbxo6EO/z+7+Nqoo85yzE3SpZHSRjRAWaYp41TucQg/EAFPm6xYIHr9etnCewx5c+MCMw
MSIgUq7gkb6VZ+ZyyKh7dA/0w2c2J8tE27bmrv2/khkeBcXVocvp8jPymvcCk8OkLDlzkJUlt0JL
6NvvNVV9m/4GquviG27+xQPPgVGX7mkSnk21hlT0UXY6hF4Y8UKJRm2NiEZFyoyAW2ZhHwahPj+W
mqAXyGAEznux3nFZjCP0zyEz6ERLK+aR/17swAwQbm7Hi9fjh1IGWS38lBko2+dbfbTbP97/WE/w
7Sc+uLrso+NlISbcCuUeslME+OqCu0rluUS53kVkPmIU1FwpTZYQ9ymGyyXNadmFKQfq83ph5Nz+
FrZWNY7pC5Sc35eyqlI0oNPTJVCbcLGjgxxyz42QN0vd42YZTSmLkDYWAxwbC5SFp5qYZrfaGu8W
FdyWNMxrcwGF/1E/NqzxsRcUvQKCfh+m5xZQ67jWOSZjokbNRDMIY2ey62xJU4GydeF8UKByNhD0
G6xt4G10S9GG/zCazvdDXNr/1Y0H8jLkMRc2UDNaWT5WTQv0WilOUg8gJpJwD3zRKsnICB+cg9xA
kk13Mg9snboNRc6SbXV9sWcuD0CQr1ByEJ5OLz96Q6H1y7q6mD1UtzHS+NV1r8Io6Gbo5ZwO1IXI
4zix4FcGNWBorLC33JbjL9rrjoVpMKK05JRmeX1b4CkqKwLzRVDMmucjkfYrexLmvDzowKoU6Wyz
slds5yZdbuoCOIvWmsAMOKFnfZfBslNnBMsGjzMLND84Dn1bCuHhJBH0uFwucnO1qvB886GSEfe/
3eq3dDGBZf8r918vaRBKwClOE1kO00HkPHK1vax9TFeGaFigUcEXFai3xY8ENHrInGRCBtXQ2cgt
L8766ZxsiSssOV5DPu1DdkemYas44LYK2At04cdA/HBLyGMa92gRj7bSGJ/0u/LZoPFnndWf7uIR
dLZTislQ9bH0WCyiVIHOhHpZ+FWcDtjj6PvQTVrx3m/v79Ub4G89y04gxhty9WoojuxQjxemmLOC
khpIJ7+npC2qY5Zp2W4U13RMjecbQdSP+8F4akNSO+6P7BjgKVAMZtxLyU1T4DjZUH90of4EU+xA
fJy2gQ/AXyDqB1I6E+vLcG62u7qRmxUfVfWMs683Dvv08PQaBmgWJ/zsJyBNgX8aUKp4sgFAqlQu
7FWnbDeVd78civWXlRP7BC+eOSM99x2r8Y1YQZ7pLZfFXPpXZkPU7bA/4/GNioi4CEh1KmE1rZLb
VYZUgPwclMtG1YKY0L+LAJ4LKP/Gptb6i6Gt++oJ0LNjbNCBqOlNmse47svUkJWw22qdQ6OhNOS8
NhMEAc7uCapc+ytfDHn4fV6fuQ0Pza6xxwic37ZYr6WOi+0QorhUgcL8NUktW1/STPlckxuM6nlq
JyRNcYHhMwYkIlboB+4i91Kcg+Gkia2zmdu3wQOVMe8JK/g+/TjfRd8Pw00Dpe77uT4myPvpSWni
0gkz3bEdpTQtPCzEQeattYf4W+aW8UGPRKSOnFmu9ORlovYaaWXNXNwNkG6uGCwb9hZI30buSul9
/6wGKKdiqJW2gCUYIMGxlgjQWZK12qqCwGqIGoQTIWOaCO7g0rvfjtEa/qYt016QH26msS24UGV6
rcBWui8YVyEEbjjIC6gNSUC0cBbQ11t2XKW2TAgACXhBffl0OaPJv/06lPb+FUKXIK+cZ/tkPru/
oNc9oJmgbvNlI9OfLt+Kp7sweteNW6aeGczNMPdEXfRzrqTEqNld3bB2f/X1obUEVrXtHKTqyiGx
YWYVIcvS++b2IlFc843JK/UUIe5I/1fJPY9JydUi2TcjoxJNIBeKGWsMuPmciEIKgR3g/dkgb2lH
GTpSrdjAKvmR4oXW+f3r8qUOPmKdHtfW40beZDwEUEAYNuGAy+gT2LvI4CQnKw45dcwmWJjNYPAE
UvEZzIZ2I/i6CnUN8DYyZ+jvfQNapaTu6w5qhlDaKLDeLAPLhl02OyjmIPjQz/VNW/1PlKp6+bTN
F6/3xXkl7CDrZVe4usG7kapqF0NpHfYtKWixh3HwT0urZMD3kRe4aKJ8Lu2ijNwOTt/iNOihz7ez
Duz/G4O9SXWxMeFLBkLbpYWnnehe9BYz+GMwrrOXmd6TvXf1NL7r5LuTyNBMeqKYYOa2Y1vjWbRM
djX2jA0WaaYtQCOCXDV6Q3etAIUAOlk1vZym2YsmCuzeRZFF63l0PgE8pqUd0/7yQg381MKa5Uph
QcvyYhnKEgOX3jz4vUmjstbfI3PsI1qtClnrIyG7XPijE5RQEviH0YrNdKm8c0A8sIJnNg5NYOxC
NmYaHyjLpwdb80TVkNhfHCzaKq35ZqXTfpljiFlczsJ14+2NXKXC9e4nKYmTR3WJaTqzBUfs0N05
/r4Le5fL44H1Q9UrZPVnZBPnDv7g+YY7k15V1ez8mMME0N0PPXDhZoq51IQWxmamD3R9+NpKBdc1
YDPc4rEFmdjLPQ2jBwYQ+pmqwCXkCYWbEsr6705QDn2+yfs47Ms8njl4iSoByg7W8dsKeYNOj34G
ip/UDBIJ093kgOWmWXgll5lGaXO3WRWx9Iea8nnIX1o8OV120cNkszTnGSxoi1QRhGCwBjdhBZeG
obaoEj6jlq8iWW2iN0j9yYWcUGzfGwsTplz1YenF7dQq5c96v1ls2OWvpIAUZQoTJbasoCPP0JjS
5Q4U1GxYe5Okpb54EjmKV3x4uN7s0hlr7755Paf3zTsPs6Io00gC3rAbWbet+mrJDudUl5/35Xxb
jzgFMNSYUJWpT9ab/ZyBGKqp5ykpBObqR91PaWEUV4V+ou4li5g/1tDYEJeL6EzPQUClJ4RwjFAN
JgFVH+vvDiJvgDcUK7FGgk8nm3GpFtwTgq+ljNF1MCb1St70V6vA4xHPua0urcB0+sN7Vxbi+pqN
LETbhuhWgUZ+wkFRnHm3P+GpA1bIhdavhMJdyjI9tSYv1x2RjoEf9eG/B9SOMBjOYid4y9lumgIt
jxXyBe5pEQJvxugFlt9xTF8tpAAMHV8onChpSldU2S/iQrgqOii57ODDeA/RVsYiP/uLXTssJV5x
RMlaYjV+8rNJAtlgXR5gNbbaXPbhHBJ+vtLr1l+1FTkzfVIXdUtMREUbod6F0BsBdoWZA0cBiBn/
YZ4fALb0Wp4HfblC8nz4K+RzFVqrvYSO4o7tRF5Yl1x8iQYuKeD/UAnolHlSVjQ/hTyWbMMV1XFp
S719B7ZpFpmqC6ZgHzwM1OBuV0UKMRdbYUFrCgvpMSbIRQeTK++c6MrUCCcFR1Y52PATDXMHtRt5
8XUQAVsYcuUnKXrSLPKKiRO2AbzsTCoUbPnbRCcf9b1ff633QLu4d/sBYmr5dWo03ytraHbjBefc
9tmVOJDcuOcwrUeKyWJlURHTtfKVcQn878JDTzdIlKjYUy8kChC0lQYCfU1TS2QnXcsVp+Z/CCMU
2k/aoNLnj7trFWmKMP7NLoSME5Ny/A9NNm67W2rVUMOw6307kY7RELv41uBNOqJDGRzggouR+Lgo
hejnhseQFrxJL5ZB3AgOd2eSl/v/j425c+cgaleupw3xUshpgppcdTiYTJdX3QoSbZRJ0xGNzAqn
EQpjm4DCqF6AGusZpzu1BOHhSx1bZx6STg4YkFoHCyVM/0Kx8FMQSsheuua6wvIkT2xGMOxQRtjk
S0T1ngGIRkHmclj57/hPNn4T6CEvOv0xXV9suWS7GlM92W58tQ4jOyXeqbOiOmfh7b3jmYdF7wCr
w4cRnhRPmsuQSjlya0LTZrkWvc0FWw65SCN+UtgEv5c5V67F/fAmoGtyo8AK6et2gt4cLwEDJErp
z+49fH+pJ+AREF5SEHdiKDJ+ZIiDR4sVz0aAkyFzFA+ys7kHtVVNkYdLqeHKjvpcATO2hK01R6wP
QSa8/i05Uy5wlyCJxobm5rUFgCNxAxFmUOj7JEDxq6eVhwwOZSozI8PIMW/2PTLiNqCTFPYX4Xcq
xr/79hYdEGrvdcaaA70qSuoEojBMUmbsSY8xN6/6/1G8wPcAz9mq7zQKHLsqUcd0Lc1qgP0rI5lO
8ixlhcjVH0H5g3aZtg9ZlVxiQiIG9TyyUur5BcgJRYTfqQTkaLsQ+YlrGZ7JX7NU/Zjy4+oI1mRV
MiNKPwRI6Xz/bV7JNASQ0awze8KI/PNRYeFwCxkVhicTFl2mw2uWQBaqlAq69Hq/KEf3zf5gB01Z
MiGWAVIRppbxNCk8dW3Xs8pqZheMnKg8ah04Zn0+AkWEcjAtCMCRAOqf3lUtKU+s9egQ3elQVihq
1LL6vvaDdKTAYg2625se0XI8MEC4s0L3ldAyTeLumWaukaiM3mKAayU6pFXcvAKbpUpn6pEvUQge
25RPZYPd93I761QJG+eRCTtKrhssc9GC9qXhf8tR+u5YKET1vbrTSBthd1KHbvhi/JrhC94YPABq
GevhRUz3iG6hceix3h+EeiWcqPpig7TvuPbldRN82etk7abGxpR46PdvCfn5ZxjdMkeXEqSBi8yw
yRIpa8lx3OT8KjEu9qYB5+w5vpMiWuofaH5IM/bAw21rUmxVvzgfyuO7WxA3z7YGqUZgaWFmh+aZ
0OdMXIkPUsOqe3ZHEVO84Y/h29oWnBQYVa38pw1wCUezMuD3NoQubDhy9LWnAOroaci32IqoQ4G8
drnydUO8Be4C60VLLWGRLrGU3yKfqeo4jnqiyYpiUSFC/Yct5qh+P38FucZho7igfFgO99JyJwOd
Id9KKEO43x7SOYQMIzGNIBlb3UStoV0yesQwoewAiuiySODQ5CwEtpCV3FHWaYRBco6zrLZbldlu
daN7IRg70/ppgzlprdIpUfD9DS58PbhcQmGPrlWk4solVxZidYODbd+IWM3GhDvtb/KBlItQlDP5
nJi/e4O+9XQOpFzfN0Fbx+N+qZYA02h79fb0Y+cQdyKFb5dQ6fPAFJpO8oT2BeZIfETgcBZO5UYD
A/EhHlKPY3A+7t5+Fow1wpl2JMTXPs9GpkxFCLznwu4CX5E1G6xyTjfWRsp190GF1wWUKXTAPMVW
nWacOVpVjjhxhQogYYtV7PBxFbqGRxS9JlJbMOLBMf/A7wceUPIcWRhc8Z2rxhSEZDsrsn3kF4Nb
qIi9hHH273HRtXJdbQMtdgscsWsCpio9IG8qvURdpshWs2xWLCqUyplDlxI6g0XJKR+IzmotuXVg
GD/tpjLfJ4MJCP/C+XqZRa6WEl5NfyuReHLaNxGJy8xx2EWwuPCvMVA85oynGa13q17dACcHoabW
axw8ynUbar6MESQYgstJGLZoRsqOxjMNz2ozr+BNAmvFSRDLyQLaLm+pswd70N1P/Q3ivua+bvmb
0dAKdzX7fPT5hlYvDWHG2mlI3FTJOrD7g7sh49YB/SRyXmgDnVf+DJPTuO62mgcusOazJN8igyJa
wGgbSYVSODr/Jq4nt/ZfpH0E7dkC5y9cORKUI8EYFNPpUbCwM9UtzdQS7ETcGLM0SbDfXD8+LvUH
Upe6EvNXsjcdvI5JvbM4JjMo26zCQ60tY8X+Hz8IiLujg+FTFycu0aZ1JwdpYEPmft61xHq5k2aW
ylr4EcEW3qRGzyCZnkyeklOL+G56p9D4d8g5YpVb8WG4ZhalFSWUt2drFFFqsMuxjtodfL6zB2D5
VrJF6GG5jMYm90WgIan50nIJ4/fkZN/IzNGAr7K6mT2/8xSCEH0Ioq6Z+sL1ov9w8IdVc99cXFZp
1D+quYTiT8O5rvBq4hq8uSR1TNOPzqMMTgEVTKXbShDtUqy4Menj50y0tmQJNi27rH3oeHWlXunK
eEAk3ZO599DHjGGE2QfOcisY+TZ/NedudWCKPk8EZPTbAkyKXCg2znd99ipmd8LoHqyMc5Bk8i8X
gpxh/aTKZH7eotbIougz+Z/093LEzy9C6YniNGg78d/TQA/ONEBpo2wRSmDovViLT24S8iVbIOS2
GIdmJPrJZNDNJWZW2ynlSPy1f5yourFrHnJYG/tK7EtCgMjVGQQeDPPYfuYkVzMQ4SyCLmi6+TG/
+X+mjWj2njVJ1jm4DY/ibMuU2bY78Ut0TW4anYb/hAu08mruSPXwi5A3balZHsZLaE96GsjxuCAb
4bT2FU3KlrJLWkMyb86obb3/S1yzqDIZN3nK0A3bHNHVQCgN8ONyP277h9GOHDS1AnLgfah01o7Q
g35WW0O8KhiZOyDQDRHM5E0+cSuJ6Vmhf0GRHnRvGKXGFrqzi74WRVkZrdwB8z705pj2WnEHlBvI
jv6Z4YmQNW73g87U9NATbsrsgASSi8vDYERgVkQ+CTJN+zbXm0zDRcdTO84jVKIEx3x40lk3aLld
QSm4FmdbV+PdohQawEkObrPGoAp55CS/oBUBZ0ZruyTAmlQAbb0Homlcqv+w6gk9Xxbb9lbo2Oud
Vxl12JyNSvGMIM0IF3MHo/65RErRrA9o1d+8HpV4KJrYQWaiVpJSA6L00GrCIaqkV6DVWInH0Ya7
Miy+UXFHerPfl67Mg0l9bMkp5s7aYs3tCkmtWSx6pxieSb2T62oO3c7F/FjHBJcyymIQ4EtgO0fb
He0lx7g00IIlVaFrJWFyIm2WjDln5RtcNvF7IlKDSaXEJs818IRTF+Yms7rlwUvTCXOmDeaRBISW
uERetWSZPXbsygNWbDv6A1jupgF+C422WUvCInt7Njea/4pOcVCwwnldH4R9vS2Jf9hqR8Y6e1Lm
EMrd6BNSy/zKrLR/orIRXg5eow/LNnpcen+T9vEeLg0mPUZ/Uno+U+xhJbkWMV7SH+kWROBiGaZo
Mk7d2TYchX5JagfOvxrFZbNzBDSoDTQLrCo+XVXXwVCtyB+pIILWYzpq5awCSVEejt9yhTDVuFAp
6uCBsHGrIjnxEId2EZ816meAc1BFle2uko3QyDCKhxkGUXAdF1f8SRQTYyh5m29BwOK4ICm2hsuI
XYUXfkL0gep5/xmUhtKl/rQgPGG3hsaNLQsQaGGOSlN8QykS8RrKSNqmFjzKScyXqxQd+1IPwO9Y
BiP03JV+JmAf0eNVf6MmUPk0IaD8GR/Q54+XXXXEva97v6iPR8bBh2dSGgsKLLfrxO76qCZH2HzG
p781vkSblPerzXVhjLfoHumHIKTGbEBQFxsjK1WLAredwTO2tfX3uTzKheeA5PEJ1ppfdzdFE/X3
1d03XdXw/KeYSukqqVDz5ZxJQLmDN+rJAXeFkYxmBu3gkEQOWBceHCAlVraMzna8IvRFSH12o6qh
u1ZTtJoUVDb1QOvQbDQoxLrnfWwiRuLIH1LsA4vn3yObOoAkFSIQolPofzuQ/061LfI1RKhwlHJ9
eNruE/cA5FKU3QRHfrhU7e9UHWXK/4pKysE/HDQZyVEMQGHKUlDVBtQynyvUMLEaeKSrUJ7dznod
SB9ICsnArNA0AwRv+UnMoA6KvRnV5maYQ6TQcESjrdK8WCQAw0dqd4510B2mHRMd/MZO2NZOTqGg
bvbg44SQPdCWbUuyZNYZQEvZLe21IiKNFe4if6wkNriXczrWIVhrNJQTMTFQQhXmgs13CQQAdzZI
ZSogCYxsUOtoJSgJUiPmCK7GRiLN7CHY+iNtWJd1NUsLLoLk8XLD/zLwFheqGha8F43y0eqKukAp
1DO/UrDEJ8Q/AX3dyGnDhTDgTAfXob3jk5DCkrt4nGPhgSVzHUZNgk0ypop11d0WTd3b0Q4qzpui
t9yqU20x6rxDf088LVVzpvVhAL5qKPmPfwvhIASeUC0U1CdfrcDvxdPtUHC3k8qzmH+1lGZMaY1i
IeXGpD4MUEk6TmuMKxRIJTKU3RDibOigbKVlwW5v61LzDmo/P20lXC1rVmSBILo7n3YZHBMwlOJw
oqE+UrGLjKYMo0ZRA9Knf3H3uh3lHa2gf+SNvEFUXR2wkS92oeNDsU+P2vYZQMpyGbKjNW3qCquh
dnk+u5AhFU/xKFw2SHkugGqdH5C+eVkJLsyaR4bLeGIqcT4RLh38JmFCJ9dnDjE9cDvqbhRDPyQ1
qYEFjiqnrg9sD7VsJijhwjsEhpPk743+jrf7xBD/IMwKLEzKoyan4PYrSFTieLCCBYi8RYR5qKTB
O6KROFIAdjDTds8gMQq71JAgVLP9XgEjyewu9E4ir5BHKvZADbDol9pDup1jvSNjYW3yWAVcgBTY
f4cLe1eTDpiAULxKzUvecplVS5mfy88l3MjO6YYkVT6RTNFp/osJj3snHRgG0dOsmkeEtKps5JgP
/7MkMifsWUrxv7+GUakaKjqHX/WgiUGhUcdQQR6ByNXrvLfLWgXpv6lirQf9jo3q53297fDVZPtm
dxL3qshy4O8N1H18U0iXZlWhotCHezjsSuT+qigxBygI2vzMdFiHYnFhjyDXlvLCII+Dc/71riYG
6Wm3gMs5eQlttc2yaCnWs8u/YfG39K4AEYp02apXQFSb6RAASiwu0boeDnseRNWJXZeAvN5l4g2A
9/nOyQy1MwDh62n0FytfccRg/s6pSVsO8jRsy14T+8ZsfGVOkCUKBxZMIbNFsB9VTfXrX0lsz8q9
r3ovnjar+IiRTuUb2e9/C6T+LPr3jFkCoZAfx8NJ9i2ERSVpmqwRhoNPwIM1lqhRLCMirimL49V1
l54nMfLGaoUXjp4uPHyEc8VGt/bNKkkrUHSJ1bXJbmxhBO3Rr6ZZCI27sdbGz/V61UsFJUnCrGyH
yVyOrp5hTg0d81ijeMjzHsexKdXlurbUo28bBZbXBAmXFk/QIxejhN24BQhzdLvtuSgQg6CSCEo7
KznJw/iG4HUgimCfmSSKMK+l7G/ziPAc/pXQObQ7LCayXiZ/OlHrnx9EokvXiqHm+/qaLgANgWDO
OvvvR/PIMeqP3jsBM3PFmhC5N7dX+E+J1gd/U4BaXVK3djvxSpCr8juGncfOrlB1Mmxz0cbxICY5
NALETjHjH0lDV2/ADG+4F7zojmNpaAp4aU4W0XWkPYdMn2RojKBKhX286Firn8pNtHqh2RygUxV+
3rID9LHu+vwpdKPtyNbo+AopRYzWkueTbGFk6f/7rZLbILF3H38TqnSvyvLWQ/GY1Q+rLBgg+737
pV0kY/hzADq3XJ+GN6PyGUY4rxGYdO8IHnJcUXwNBrdya6ERymlpRlZNQR42KpQ7pcft0aRikMdu
iUsNKt/Dbg0+/Ja40BY8xXhsl7U45sb2PvJno5GOTGxAUOIMKCcOCNrCNbDowfYQJ7sTvz6/39Mf
+d3SvXXsDI2dJB2hqOBfE3/WIxn6H9hNnR6oQAzyEGXNPKrIUKbdjdyF2q0zldoIWvqnwuNcO4Q8
oj5KC0Q7K+MGPms6iyc/P4qWf3iimGA4YBrKFqd0c/pljTRaaNkxC+xABXM2ZONnGXY5DygNxFWP
VkCb0+kw78WvaHPNwnmmAZPlS7bYWW0YXqkl+3Oo+zDFWgMWYxV0/zHx3ajqQKgmFowT9UewP79N
z1pxjaEaS6jj68eDe+drRKdqxAqYEQeI34FTpTUR/Nn9wyxCx/E1EsdWNpMoOqGl+AFfGi2L/IaG
WCkhIbzHWehzxWlg3Cvf9KPNLJ1yiaJ6glKXeq9f92jO4LetN03qsDWtk72M6o4ox0AseO2C4heK
mQ1CtMS9MzuvCevtEoJXdzy5I9zlJIou5T7lQCZqYO9R4Q/V4SKCx+2tshXBjuuNIu+idtcvz26F
niJ/cXVHFO2aIhdxleJzP/bNwcfHZVNylw6T4pbxLlcOht6cVQQ3WvZoy6oPwA5Hjs654AsuBA4q
60+ceYXayl6sQ1Nhyosu1X0h0y9sAsIn31SI9rVDstGlahm7eDP44o3y34Zlb4nFYjG89xuSNmTT
T055gcLAb4Om22V6ZTBuoX9VMN2fVh7/RJtJFBAQWcOsRvC6LdP800ARRwdkFtJeBVxM9an8zcrF
zQSawwPgmJfP465LkR3pE90Ks1X4HlaTxGGQ5rE4QM9c6I8qXAy2fsYVaWdQAKBR09LPls1QLuq1
NTAdiD/Tf2+1kJIPdAkrPnzaqJE7JBCaj5jhw1w3k0ozHdet41vcwJxmvp4BsdczAkKafvSX5gDa
W7S+YVYIgoX88nixAZtCN4DhisE3qkJvP49WFlCTjh0rfIp5DGj1Tpzv2N/2Cn7E575lx8ZvXo8h
Ox6M8SxSr6YB8n7wlxVdXoJewu6oL3SjbR2nTLy6UIuukI1rWxkBVRvn5ve9Jv0R7E9r0WdhV4KY
Pr3LCNFI67YyqAsL1Is5GojlF/9S1yM5Kal7dm2G8DfcV0NarGssnXLKu+OBzMPwSHQ7ngzEAjjY
sDMX4YsLFxqdWfE01LPtXVVXZs0mbe3P1Lcvv2K7aD2LSH6IWyUL9T08eVyukZpDEmNl+yd+oJxI
m2lxlF4J4/PaKYqgw0n8ToTJXwNfB0akTybsN6awMHJvcGyj3vf1lPPbLagA+mpjgCLMhLf/rjRy
hvam49aOLvYcQ3yB4s1mdswepFeRiA3baRJ9OcVdXPA9jZSgI4AkH0P45F3yezbiRE/CzOW+xsiK
HCqojn9lhXz7E0dfQKwV544oZT8Mvyz6Qltpq57UREUP1hKG4bBuAyqvApEgl2B76BHEHODB7LcE
yYAlazJMnkRMbVJHXqAE/AaryU/EVSJvFNIX+lX30hL0uBByJFNK1z8RaSnZtiSgiK0Ckn+9TfJ5
elx32H+6iSRoIT3OJDwhJnX5SkrXU4v2bEIn2DCxa201oUZLE8kD1RLIILjVPv29/2F0k4vXNitS
XYPAvQfJwmscY7efaNgpzna5C/Fi+0NcQ7L20U2u2RdmxEGtoCoZHT8ZxR3lLkLZx1gPPrLfYmYZ
cBnyEeOgwX3KJe1VNpfW00SNr4aFHrWzuUS6uaOwuFmIwQQw99r7ue8+hkHbkJP/7Kb2xcO+pGle
frC4FqszP0/T26OHRLGkwb0BJUFPu4lpRQyCp5UCXvsuCR4ejtb/z9pKuP0le/6RLMrVgdp1jWRO
CVNkRQeBnok+17ZS0BGatp0UPSc+jAATbnUXSxkf7myicO3Qx8MI/t+0p2iAlcV0a5gZaP9Z8R2+
fX2BaqDkVeMCeRBc3y+dPfOiWz6TVub667sqrNXmlbOuOElDniqYG++U4RrMcV0eVVE1pP5QqefO
KTL5sUzUI32VxjIp7PljoeiKSpnKOwAYogtxl+34j0ZbbDt24WWqWEkFwBjt2iibni5SDdbvjXzd
CuUyM23Pl4S6OtS5aL75sS89CukDt5joHEUQ5oTT7IOMixtAF0cWn8XxTb1pACkoD2+swSPEUvb7
pSpio01q/BiPxkk0ogQhjb/seioatnjWaatj2v8RtDe9U0AeK/QXiz9LDZNdhDIwTQ+32FtCNsNo
h0TGD1s9F1AWj9f6xoXqz72rZdFaucGHHKt0dd5BG8rU4RGHrjR3ejD/fhpQ6+1hZWg5oAcTcP2a
x4Dng8HeOChd0oX8Gkbo7ZFp4uI6/Nz0HfpUmNrxrjPEnOkfmAHVqECMEflOXtiBktKbtX2s0QXQ
bFQWlpa3tAnzDV9MVBUvVv4IBRXidp8b7fjj7f1we32iKKMff93PFVUMzl5/dowt3Q8oOKx2gKF+
5nByiKD3hJjpCaEilab58BI2+LFWbdS/RQvmz75uvSbnsi1CtsbVK46YWAJg5qjNRFbBzzIpGpOG
zu7pDOa6Fo3KkSF2o/FBZKKy/CtwmBMHRucOsJZqH4rrRjXCBUPnw1BJS//lI3J4TUg3urlsnOXq
1Oe4UnK68pI7yFMbzBjWZAyjhDZSUy4cY5E7a5zYBsqrUF8TdjABE4XREI2dXkuddltRl33K+vJq
iS2LQVasXgsboh/WAJeG3BqiiHgnWpsBR26yXV3ESFCjU+S8cXp3kOPIWWg/wxCoeoDf2KEAyGyG
ejSMxgao+Cdt6hb+ceWrLvaEcqz6Z9hM2OXP8NnBpfBGPbo7KO+EBDfYU6TG0d2Roi2pKtldGyew
k/GJjsYFG07dG5JjJb+h/Dl7UnCqfayzBQ6JVqZAVmx0ECh570pvDKOrBIDcwZbubfeTe5Fu6QHT
gMaMHQcVGlHiMadeuUB8KGYdfKTcHFxwo+kqqUTtxHnlFk2CAPHr9S9u1Yhp3YKo0XjDex991yAC
9D8nWbjImh0X22e2rPhR2kTuCbhQCekVodqndP73RVG+SPxJhmhqV3wN601obB9eGNav12k04O8h
MUH54sjMtr23Yo97S5r6zidElGL17RdXJlqkSJC7CMghC9GolxfVNZ1td0Fs3oEwjBbe5XOCRuDv
6K2NHlVEYtZgHL+VK8vBZnjlvH+3urOBxqgD8fnZpx5QnfE7MO8EEjphGd21gzWLIZtWRR1/8j/I
N+jj2QfdBvymJbbXZVnvxsqV0T3icBaq1tMCG1f+y49Ewboe5NfqxbEMWB+K4krt7ZeBcjA3ytKH
+F2OG2sdbeX28+XZejx7NHwXuG/6e5kWx1iWQ1LLV44Xg5xST16f2vzs4GHu0QSNAMkivrZmREuM
9uY2/c8y+01yzftwuL+tTmeB+Ljigtww+RO+kA+Kz3TAJINctqyMNNlkBrT83JLRxe41nVx15x8U
YmOdGu5GUsgFfhvusAko1bTnUyd/FljmQ/ICMWSTMOAcXcmppoHRFGS1merxY1I/LrzsMBzyv873
AiAkf5q4pfdZ/GjCgHmraI2kFqrpFZs7dpB3fL3ZBt3IoiuMVg5fJcPj1ux5xwuCPVERxdurOIJD
cm8bFuZd2dQXVLt6G1p5Eb4cJEmr25jlGA2NqhmfM3GnQXP2Q70H/YCfUQaZGUd6n5zrpmYEc1Md
l6eiVgK9qG6FvHlo2U3D8owZlyVtbibKMNmg1J+FfUuly9T0bjTtm5DxMNAgPoqHj4qtKt4OMZkt
KCt3h+bMGJoVYBUxTOvpNZap5xlset89kcacaAJmuRKzR8nBP86i3/v2nljKS87OtcUBx7NPBbX8
amfgfjr8wQ5uf3PTcel6xQKjX+290QLkAoQ74lMUcEtIyseLwrjKechp1t62wocIWBtEswJJwTQv
RcH0sb1bwwI177fEUg9xt2Suo7CWJsyFr0MO8g2MskDtYQpM4XmsmqU19PCd/ex4hLd0QxEREivy
JNLcjLi2w9VAHjhjDD7SwlA3tES9HZTJXJyxlXMSRFDK+pWoztav3y40joXhssNMg/Plrguv6qMF
i8aTxdAjn/L+heErzwjJvVxNCNku/f4d9ar5H49amMzodtH3f0LMq1fGoJyuP9fGndr+h6mInhgN
GZssyUQI6rzFTpwJfYzI/ycythhWdL2aLJhvJJtil4SS6LgQ/iOhXSIMWUme/Xgd3YEXBL9TWYd1
CECudGav51LceSNLOD9h9KnG0TEtNzgm/Z7P0Ful5PUUeq9y+VW1y5MNPRnyyQDGGvfYkvn35j2E
JV2QrCMCiKfS5HoKgXCbygJDu9eFeej29QdRxJG3PLCVvC+MCs/7C/e4EVAQkrVvsP1qat5kv7WX
I0fYVwvn1cBFmtYUoXDWyx9NesRes3fQ305tW6N/HM0pNag5mN+fEZgUljdaWS92IqkzXzHZR87g
EFZDKiRzA9XT5je81U4j8S11Et4mUpNzw7SxFjELjZburJAwvBvk2xoClppy4YaIqqxXOdGJA1yw
auZEB2fL7d0zUPJEYfqQI0pKoRcr7OuHyyzvQrgsE/XqBVUjw7G9esIn9L278YzuTWkMLGKXqpYv
1i8Py+oGGgR3Zfqk/bnGEpoltYyWLaQ3VWajEtRLvWlUd2WqkA54yxOPTLdoQHMPGdJL1toyc+sI
of6IwC/jm3mrtVe+Flr48vv+4ya15ITjSvXL+btYJkM6MmvSNdXOQ7xQLkkzK1aWzXtZlRwWSOh1
xpDchhpSRqVdcN/RAt0mWwQxpm/EJT2s88SUcH9Zbvb7l0z4jWyMv9E/eYTcvol+VKDT8RPvhTAG
+qMm19MoVhLe8/qBLJy5Bq7TfIsX9IF9cVhYa2y+HU0WJxsDe8mrCMf0CEPfUtnyXpvSolq1787I
Gq2Uta4RPZB4YsEx8E++xl1WxUcRrOPUKpvmD5JyoC39vrWApEVWttbiKrbuvgWdt152rN3NwW4V
NVz7lLKgkgqO2aknUuw457+eJGEX/fkJfzYzBqexJJOe38VK3otaeoehlVn3hUaNRNVJUUbS74Ew
WQfonCZhwJ3cVyUUmJC3Ik8+IqGFwqxPLeeGcnSzvigQKpr87EEuLT3XhZqOiO8duTyLd70MIZUi
UaM+jb9JmeF42v25KTkP5ZJP0TtYy7Xh7dBZUqO17oCIudyYn09AWCHiUuYaWKw0vsexuQLcqvQm
pEBCMabAUxzxvtbna5X4fJe1f5FNbVQobvkmDLC0wuhwDaLCvf712UjzQrfYF7YQHtCuHQVyQ9iI
NQ9GAIo5CL0ycRPPwiBQZrY13IYCsGujnIdJqZd0MLhIHdrRnOgIBRGLzmUOo44LZ0MsKdUUeePG
sdQk5Sj2xSs87IJB+2mrM58dwqMdjpQpNHDpbjvdnmuwiU546yksyyEG9PAljWdSnQFBRTISL6bj
RaRY5ohfBSTJXveEih7AMhT4/aWYlk+jnaiTaNS/ka1ELbfci6hLv2neyzxVOw11sgbGhoXtTWgk
6jzNxjeG++IrWkPWoEAJEoX5Ny1IFHvjkI5/DFDsYUmGrnC7pyIpZBpXVo6JWs18CO6zDhVBQP2N
dviSpgSJ54nKaxWZIlQEQoTzhGa3mIm4ZkKd96CW+LthYFgv6UjTN75vbkoNAB9jkTHygf7qERIb
IYv8z/jdiS8plbDKgyU1g4v15AZsDXOr29qalxv3FQV91F6QOz310jYTsgVT0Qw9yrCX3ZHO1XUJ
DMgclviHFbjmGsGOlOAyKOC3VfCQLaDECdAqTR0Uzs8TDZr44QWpP2foVSj+MQ7owxpuEd98IGAj
hX47TKxgycoTD7LLmjf/3uQ+QyJN8TKpmaCFd8WBCRfxgigF6gx18sKDfGasmLLMv4CK8+sWtlYH
SmH/D+c7L/prcYqUQwx3FYd2WwsUrJDtOFLfk3vn4yW7NYJPGVA/TAjs8Lb5pjBnWNCXrLV9FNrP
fxnEJtyDzKIfSO6q0wYHLPXw+fQnYjJUs74mGz18UjtF8K3VJ7aO71P3Ieq2eJidpC8sXCpKqaKm
OKq2lgdb4fEg1NeErFXOOifBS6Z5teIb69uykN3ZimP0rMLFp7mFYMJxR27Tgp/gnx3y5slrCDm5
nCcXIjLMUji0uDAYSTf11Idad5XtxtUpisggA/RuueGLNVhVvYBDhct14LTwTSyuPmQ7lhbZ3Avw
iIJIR4wI8pzmvvqadp1eTNZiDJ1XSsaFwFWHbslTJxp36jFWsokN5VTVbEV5a6DylJp1E1mwurUX
h/+m4c8OzTg6DpXfsHdYWCrWF03920Ps7VKDNWaznwxlH4XemZrApR3TuUjc8jE3H932SjM+GrCr
lOMdQ0Su9STDd0DA1OVmL1EiZMGS90JG79Z+nnNApWxVA5nxfxK9nOGoZXFZwgOO2r2o/zNC6jIU
C7qXnmVVoUPdysMnmLgBVZdpCwq2IbIPeug8GBCqzeu4NUvWbTQMnl3oC4mBcdxfEgAkQFmWzwlF
U8/C+wIkfJI2FwTOYOx1yBjkOVNGD7+jTM4o3mzkSdPpZKaNbnkQy7UOZxWj6MhQqg0bXICDSbOf
eZXZeAjYwnL/0piARo8NASiVPiMjPl53wfPrFESA551s0k15/QIjrE/HwTLYUi64H+6uADNRVcAZ
oKmvO6crwn2nth5yNa3aTudu/lshy+rC//6h01DX4vXgg9IVK+v0QCHF1YzmPYTE8+LMdy92WKkJ
IOjG4bKEQQfQrOOibJIIKk6Cb6h3PTWKcdpwZqf9ycPAmARG6xnyeM6eMsEEQ0RhxRCiDHmYK4RH
hnnZldTQhXNiQaPfPHhYllVs4ct4IPNZ8WGy1NFNhrpgRZQ0qqaDJWf3sPo5h0s5ZzUZVclL+5oz
yEI3wn+s0nbuuGN/Uct731xs0FTct28TrvA+/TCRYcHbpT7l3ravPWOBEIeov5CLWh7+2vLIxO11
mQWjsJ5KmCtPG0D4DWmBTqomSUeIf7Ug2izn72PEmL7atgwOFfXNqbidru2ujpayZqzTu5mcq2mv
lnGn7WXe0hw6oDUJorMWnKUcjyFEL1BOYti9F9zcwcxXKMwk+jAJSoBQO4X60oSMlpOg1AOH/37r
3VRqWMBm68ar3o0/7nUMm3bLhjigClnlJeJIxTO1mAQ/TUYqCxuTJjnE/n4coUlVKy664a5k9Gmf
pDuBk4rVDYlYpO7J7PKxJyMqucM1VlVI1BNbzrYG/s4X69mKFWMStBTORAkJmBy5bRgMtdOFHL4O
v+75yJG1qDdHXbqe8Lu8xFK7E4DroVVoRyZtT0bDwsHJ7+34Yli4VRwRSb+28ZCu9XiL+C/qQDb0
9+Vrbrkln1NOUz78mzwThPM46Y2vr5BhlNpilPoDml49gaRszouj+NoROKxq/2NNuZplMiXui+h6
Jvz9vy5IiX7wN7pFVSsyooPRL7L51kpgQqEEmCD+tpMct9LLL+XLuy3wBMRHO3FDqr8YbDOWc5Az
qjrNnRzETVqIlksuo2YwlyUWVEeK6urMos9zqNjget/rFNZfpyodfHVVRrZGrOKHQbracn9+/2oO
0qlaLwhbUSZUzOfM6RKD8Fhv0vHmKAXuNXqmPtVrJAUU5CUUDw/zQHKlBVF3/LvVdJ0+LJcVMO0C
iGQi0rIa5f6OVMIF6S4Cl/Ug3bXFf71h/wH+hhj+Jx3YbD4ZDtR4Gb9w80tADGL1+/Kq1llscS+o
KgbRurHU/FWwz1dcglBmUb1xLD28FJhCDl5cRvOulaj4u4lUfJz7NJGO2AtYNZOGHDPk/ET5XIwY
iHjMr90LKFPBoGJ/FMNRLK5hf92BgojaD0neZOlQZ5yFCdhrY0iG6ylr0TKUKFjJK3STRdhdRMnX
uwo4uJuOHnDdr0Lpv5e3G4Q9cgyhJ+A2XKGO+V8izZbUG9GUlDNbPZoFnpxH8lS5e+SSLZRweBKE
wSF41H42F8yc6C1wR1fT/1CsjhpQk1uilYKUqCV8oP7CLLIlSrrbvpHYyg0drr7PDLAGH+rE8SoI
pWDqwzkzV33mQu2FKnka03Xls1OBbsPMVPgPC+SjCZX1fNW60n9SFI8B/qZZT3l97vF0ri3jyn6N
k7DNvO/bH9tXb+M+iubpQnC+92jeSPUOOYJROk/O1x+1wwEh0C8UtPRUViieqWysLNi4a3Ma8/pp
4ABAskWRXXIOszsaKmPfdfLLiWnSanLZS56rGg6lGCp6NeRuGJu9M4snUx6pSf5b6ZKzauuQJPQf
ubHEBJAjAKD+o8SPXDtj/v+QonvMKE6y2EAOU4UYXJ522/mO+mmsaTukndphmOCxiJ6eg7V9E+FS
tQKyFnKn/ECKs1yD/nb23OnjTTNzfGSDOUoNAAyROaM0BfFn62/HWdEOIHu7ADV0OJAhDe9y7NP+
sk7g3qzJS2hAwaUX2dh0B4HfXv2x+zkgyhvDq3CZ9GpjWaXojGFjIy4AQulgx/hOsi84CP0TVfGg
LsPvnS1rUORnaJ3fI4lZqFN5BiW2BwlGUDniamxGJcrEFGjduQYKH+fIntLtXicIEi8MAiaI9VEK
p186Qtypbox47+I33r/EuZjsDvi+m/SHfxqmNLhRXiluRpW0SzJXvDg2Sb5VjMGsVKGpslGDz6dT
P6yDWrH6mXWywpPeP9Fcm6T5H1UQcNnvoOa1ZeC89D6tUFh3cmRLu1ectK+4PXiEwqfA3fyfLldN
SjfoUQn5LY06/RBGdrkFY9mTfBKIuf43LcBbxfAn0LAD2TuS8hXexCMbGvbgLYtFOfwVFNJejxI/
kcfuVPO+5k/9o58Z9DKDtxPYa5xiwjmq1KF9/dtmcBSP1RovqqJ8kOF3eXBRVI0tcqFQiYLM43c1
EdzAmp5DFHtaDiaMY7GCTuTYjKb3plZ6Or3GKL08IwczMPanYtXdm9JAAJSeohn+Y4jePYdzZjv9
bQEzgysvEetgmdQtc4wCgGANQ5mkLsP06urMBo/9C6fV440uj+sBXmLmkY+SwDsRq9LY+sW8sVeP
JpabNVm1Oks4pfOJUagdK9iZDMw2yYwsaLDmnnXsBmms5pK2KPs5tIIktRMMqWEd2MCywVPa2Bem
ZcIK67EpHflaY+xwkyfjHn/J6IYLgmX5IVNrWPyf6aw65ZUXq0gVioOVY/44scfZV5mjTJHtL3P4
+hKuG3xyXyKwOayNQhrLoIHWr90NONa/1QrJQLJkqhb4I/AN1edKkBlT0kAfkx7YnD0SqCyqO3zX
xmt5Fi7ZwRy4tjNks3ubwArYdfFT/LC/nAY46phmW+3xDOay9YhKFoZp156NNFVrKHHZpGSHRfj/
ofsTTlYiy442hMOgLRSRgtU1fCTN8x0NZLnYRnIsX6IaYLynIqeC62aDVa04PPW529Yf16ZAQ2Lv
A0DuCC+W2AuX9RYA95vkt7FgG5d5gaEGImgFZOUNvjE4E2vf1JJtjhu/bAZ35u3xgdLw1p4j6pm0
c26Wj3a8GRM0kv6aD16LdJ6+gvZcdPxLczviY9Ux3ByBMO5nFtYAyJQrOinLnqKJ3/7QBMzvi2CM
VZMDrm3zBKnbimQG3/vPELmctYU6kT51WE3T/hIOOAQ3KQFSKKL0gL7T+anQdk/umuxUKfr5Gcke
oFnyk5Yjdughr9+6WlYzLMwbYYN8tOwPePFJcsDv12sxwDbKiWWCu64P9WxofcwBLNOozNuTnt9I
33w6ic4WmKXWVTEpNj0hTu8PugyPzLrFeufopio5PI1Am3+b6V4+ccXhlcn3FEhDnYbAWsHiRCh1
kwdCsCaCsmLZQ5njzLnIkgm0C4sAOh0lcxhWbJpg5Qjki31ycOytmhZQoadeM+XkrFPuxcsDYCbU
3vNc9pFuPQkAsDRhZIH6sb8oPjKUFWUyi23gVFCblEfVpzPzBqurTUtMDSLWDtvyK0/WTDwOcMzS
p6QBs9jWfekhuUnMcGvhVH0Ez4/GKKT0i3LhyRTGh+En4GwUtF7J1jRR85+9WDrFIy14Z8AZaCYR
Xo/uCPn+jPaX5u4Lz99PEMX74JtKostjyNe3AJg7GAfQPf2FcFCX2gBHZdSQT6XgV5kDCwD8Jb5y
lEyle0l6XRHpqZS5iuhZduuG3GxmFbXdG49Ogq0MqUrHH3jRoVQDPntbD26WWx4a6O/5tzqZmz3A
q8IFlODSrbAnfDljTVhZ7KOP64Extc+Yznlz0rw6MnGzINlW822B48kpuYEtWmeYFlaANUImOrt+
aET67JTWDsvm8y7GLP22hXGSZhJZ8Bm6X+yTmvN2J9raWWJfJuYEqgEuzSfwbDFETUO69BWgbCRj
UjCHnpLFZSh1solSEZRZp65nXMGEuo5EJNPwnLesuNLHs7i41NvMQEosB4VBxE/t0XYfepCrapv6
Km85xoOqexmVsfUdewkdp/oVDdEkgTjR+n0o2N/ehYL2HBTUWwb1M9P9bNVLp6ntaL0W7fjr6qFE
6KNZy12kiwzYdHVO+UNpBabXA0PrxqV7YY3yX6Oy333opsCXIxRH/jog/+6U5EBtJ7PrWXvA5/Gm
g7nwqJUnlMv29etpv8OQEXFGsg+rxlpTN+cqJRKFjiNQTOCKQGt81HCoaexs2D6PDWoF01VjAf9a
Lwe4AaZdAlskbP9Ij/sn3NsoNWByCVr+Srj3QCSerJl2B8i9jC3WCx8HmzfYPQAaT0AxFft9RFuO
pM2JqGVmP4bMV1UtJrF5HlIUMcJhsaJXg05QZLu+ZLy8hMFyps0q3X6cQ+jsyKyTe2wgvRWxyiBC
e8Lem4rkVWYvjY3BNlfDRMI40qnbXuQIQZFT+Bf2DLBqEA0uAnsFAjgojxkDTrICN4Tg9Pr1AFOU
WPCho/ZdiRF5OtfuBcx+ks28t1MW513QA+iGyJ981pEpWulYT2arb39sEqntO+dwPv14QefgDAMY
nVo447lqXniLhVqWeBQ3hXB3mQ8OUoogMHp81F7r3BUI1U+EPYJRJtXXOTwE/3wcUvVK681PwAJ4
R+X3s6ZolwwedDr0FNSDg3emUoGvB/eOZ26AMBdughrwO82Ef6XiPh+EyZavbmiyRZczcLWiXs72
u/vKvS66ncOHX9n/R2puCLrMtKXyONhFpjJhqDjExMXXi/9B0DGIDPGdsXe0jnBG4gf5E47fxKJI
UaERBMKLf6T2VadOy5aIRi9U5gv6ptWMo6CqxXJmZA881MDF8j9pGPXW+5jqVL0bWe30SyNjI9qE
TMg3LnUOyYqp3qa+ACr3uYuK3CbXwU8W+RIbt5Xodh1KhQixhXd49xkA+orKGjE9gQA7UjtnQ+xw
IcX4PVLbBTR8esVhuDi8dU7XoWWvxQYhkJsyuUzHw6lwp2tV/yjioZ1L4+8bGMfo+hvOxeO0cq/c
PP43XzvDLGiJ9jp+IHc1+60bXKVB4qeUpwMW7gQojhJsQ07k5ZyxRntjVHRoBEZj6vxeHk1FGL61
DZwdO24UAAnb9FAisoxfG3mOYwLDwPf6o8SjskpI7DRzkiSOaTkOlubVikuox8FtsM/s5VqE0m0G
iJBRyRq8VEFXShpREkTjWIk8dA0aFFUFQ3KGPjGoDQxOSybQp/9rz+pHOIkF/NXpHMBe378W8mXe
64QJL4c3kMnjEJ6X8g8ngolzOh9VOT7ptq50oYdGuALkkIVXvAUjVFMYfHwPdRd/bps8RsWHShWQ
OH5ngQmh+NlJ6krR64M9JZCtG4zj5H4IH/QENgRYRFNlm9NBK5HFdTPtAOOG0QL79JS15MDish0c
MDuNDkGaO3e9XPwbZtmhWNfIGQ+KeLOIr37P7EZO6EDubBD0fengPcJXKGBcgr8MK/Ku87TWTVet
ddWeYY46IZ5NnM9bqvTC8ypDoQAOULVzE6dhw/rKtCL/UNvhvigyrOUpretxCu1hmr8sCVFYFG7R
WS5lGD9RHtOT6sJBTH/QHgoUYZ//H+Yl4Ml7to/ZJU1YEfH9PiFF9ZH6RumhhFnVK5L4z+EaZb/1
HEkkUUjmvf2G6X3ZDxmOVG+12zdmO33EX67SlUYppHWoKfX4rshOwN0NJNkGLMg7VcLEp0vCYi7Y
QQawZUHLJZ6SXfv2fmSew33x7OdSvRO//42W/prwY+/GHGrLtXm9ojCp5QRYm/kSS/wAsVpfRish
Q+nkbWTaDUM7htsXzrq/gPC0H6RHKFbitNf89NL7fn4DIJ8SLVj32J67cfK5qPsXu0l1/BvoY+KU
vL6k09gyDBjk0rIEMPVdNIgLSCaItkWQgEp3zRKPcFbu+B1/plgDJfbi7d0smujt+B5TcXw3TUVK
nq5R2QgpfG8eakxrT6fOksjrODA6pRaKSaOLXsqL5HIObyBfo4PRVJ3u/tW449QNsTOyKpIV5Az2
l+cTa5cwq2g6vACKtd2ttT1y1XK0ndmyovwvDExivrX3A4y+FyD9o2uAZA7onouaee2cJBscpSPE
GrZyeeWOC+MaY/rFf9uFojlQJ5kuJ+E1aV06b9UoLmtODSSI1d7BWdN0RU67hJW13gpXiWnsSPLt
CbEce8rDxYpMfQeyJbX5DEMxYtA/Du+tY59O041wR7whUT0b9n+Z5Y36xsZ4MRWSRds1nCXVbXrR
kQUcZp/T7yQPDwP9HB7qTcusa/Lz6gLET3ZWIUC/6UGEhuDTSevBjtBF8P+bqp2BWVPnxb5OdL88
2wIUvFV/D6YVgRXg5lGAnB8cs8CQ7mOUSeOXB/BMOfrL8TxjZa5o6fbQqL5+RNp8KfkszWe/3lFI
robpoP3cHVruLov2U30Tf89YvoDV+t1VwQn4gOLy7eOuMfwRe2xcvZ7leQ+pgliauZR9xgiwIy29
MSNnJtQUsL3jHk0guORNC4u7GeFurSV99tIY52cNlsRPRR6nJQESSbkWrdhGcJMzvS8zKGpI+bp6
pfiBB7fxqGov6wDzxaMrk7EcTGvdxTikVO8sPYA6JxhpNaUfTwnxyFlOfsdwU1dTSS2PVEYzUemw
WaHU6vyj2H9rk/5S+XdrVep+3BrtwMdTMrBFrbWpG/n40/VMKugWTeVnrb4PSlvhf74prj9k3h3+
+7EumaTwnTRG5MZzzl2qpg2ULLBDIeF/gGjZPlw0r3QxCwDoLdf5AEwLQBu19rlP//lPM2Ws2KsN
b7bKufKugIcVQuCDbK0NNgJwuHIb+ZR+05v0yupLmqLxYG7z13RSCf02wj1/zxMU+QseewKkJYhR
jSBm5jEARo8EdwAXb6CKynrV9n/woHQ0GOITXC/aeZv06sHJtGQRmhAXsLc1EgPxA84JwI+h64bQ
HWeTI3FUYqFdcJVjpj8LFYpSoLYN/8ZnVk1/CW2VwuaVOC8Ky+vq18YHrm7ijPteeWNZCbJMuhiz
K1VO+AfHyv44tDJNgCRaLmCn3ZON9Q794bzm6QAa3Bx3owfzCv0yD8+/sshOqNyOkt/IDeVIDsmI
yuFBpCxfTHpPiO9eAj98m9+kjhGw0I4QPmEvheFBl/sfSvQx0o+l03my8f2TsRswjDoCC3HMyElI
u6wnjkTotu7znh1nLw5E7FqNtbNkQ1ADrcGn/e8xWB3HexyEwEG7YNHIKLgh+62djokSKx3UzH28
DSIAKL1d3B7yCPqvkyr8eKxOppwR7TMJ3GOWuHROzgawr030RTHKR9kfoPp1mE9pxYtZbxtCcNAX
3D+I36NyT06aAIPRRNxDt0bhc2T6kJvzSrOXtYos9epew4LYRhuyAqL/BZCgNA1Odzr3dmptvw27
vFJX9HFZd0SMrYD1XEjg1d1jN7Q+Dat8g6xYRxiTk6xm/vKKuznkiPqHu0YVT4HlylQX94ycgNCr
rduOQeF22R+Rid+3RgNhQZ1vAT5DMMMKBYyNeW4n0m4eWaOzUl4f3H7wn4o9rslU137W4a2K5uFT
AsIAqJAYFlToa5a5+dBegPgC12UN1mRKDlVhx+w7+EOuf6lQWAY1BPonwPvQquLqv2sh2NcZ38jt
1Li7cOMOGCEUCFnLgp11MPbrrU8x8+o4bzKJuFzDYPYD0RlJOnvvrJ8MO9bFRo2yO6fUL3iaRfcS
KyDXnHrHH23/QRt7/tLWykw09/hG2qSoAnM5+/NTovUHjPy93uVn330NnfYtC++5AyZPtBBSVbXd
EOakkwW4kESe3m9cMDRl+ri212d3MzidE3FrP/Zk04LbSupagdszaQxC7vDHLav5yMxUm6RoQgIM
IcducBqvs1J1V8XGOvnTeqTZXbFIA/Kljl3NHBzTQST9v3FxrE3rXAYCDhBoSB60jw3oxWns95vh
Q06lkkN2YCE2rO1nQJLsAdzH0wglH3hmI6rkKdv1+IJSQ9q/XeVEzmNVqkYy0cHdI532+94uPtgo
CGmPnHRTjwIMw3pamVfUtfJZBJSWDae57n2Ld2amtnxA4gx8DmeVeRfayog9O2WOsbHqSQ8zRqlP
1YshuFupAkzRc1jHJcU/l3J2x2Zg0XVZ/IcmsU0Moer1MgGbGzYzDJ2GOmbis149Qb2UhLhZ7yhD
R1bbaDFlu54pv8earvo0xyCoiIJ3Trd1cs97KlQPNoPkpvT76fzICCMKF+jpSjfoAWCpGMHVc/Hn
5Iwl7V8nqPHlBhtv0vxg+A/msZagRkH3m3qV0AYFFnjXICQPY5/o7fsbodjisQPfqQNNTyYB1tqq
pERGl2wgkSbE1gNt8IZn17Kx5NcmdvD+v9lUL4QWW8ntx51GcL2d5unxmCMaz+5ju63W3BfQzn1G
48XJZBuo4Dz1YGP9lKnDzM/Rkv4N1IhqDuU3Pi8UL7HjTd3p2AX1msQfzSwJP1ISomEYaWbxoNjl
CwIhh+46JGAR8Mn+UIToof8G+tna+fwh9YkCip9tfnnCUwekrW9RLR80PxHDRI3EqHuaMe4gwDcz
O32RwE4YYnAZmAgzR0A1KOvdjKuOKPhdtfvWK8it9y/virsvuInD8JT+Jfe3aokIwaV9WKx+9U5z
5LQlO4ppqLhkMn5qs4YLHfeSXgI3kdoKvTWE7B7/M3e5U2G80mIvqYUrwmUg2G8zauuKNZBQ+Zhp
Y+5Cf2UhxRUccFP+ys+txSocFW2avZRPa3dqClX0ddRHGu2gWp5XAnK3AYcFabNZ5YYCrPdJzXLH
/t8mhRe119zKVqGzEb9cIF5b39jBuK+LVMRThBpDs7ggHpIiHvdmJ7tyE6mdpOD+B/S00VMBlydj
d0qpaBKsLNnxTKlnWEHVIN8aXk+15S+M/yAmbHGDCWKARwZ6PuF7lyH71w8JGnhNprXkuHJ1XEyw
oARImc6JCm4MYr9L4y0t5adTT3k4M/lTRyXk/qvVO1PVwKEr2T2EILsS7dNhIhU6Q7pyWnqE2coX
nFy469L36GSa+4Z+M8lUtZV9KRmllS2GiK72nDQuyYg3gFZYqj1pCBL8AbgGQc8RDQ/z6fmNHyIc
Qem8nxx2WWDtfUcTBNemvUXhbklvKmIhPmuXOBy0n7J4NOF04QbNkk/NLoQOyHNAv7kYrIpb/hbs
wIgPYQ+KJ5+fgZ9rR1RkZ8onAkBYPThpk/20DlMVzITIsVZzJalipBWimsOW/7eS+t4gt+uHY1A4
dcIvGRgPNmyeYQZ239x2Ll2sVUTtMTKi6Md1wq8FJ7Iu4jm8lCJFT7mQl/MQ5Yzq8VxLlz6AAOob
GXqWXNVaJL9SytiDN2+M+L6CgOM1B7WK77redL8X3NwSpJMsiezoTneWuQZ3GHzbpmCZ95YhAhXE
IAskGgC1NGB8z/i5fW0/HeNjU/e+ofh/iuuOMhbpg6TqZ1tS6mkZy5k2ehKJtFewN76Y//nm8+vU
vXz5VFL2XaCRRosIjqWMNiahfyrkjOXavemAGZhpDLkdRjmMKpX1Du23kmvgmNnOCAdyqXMDpunr
PseJSs5muALjYHspgdeb9rwwms+oIXdBiMiuNfqc84W/GWT6wlccwH/DHXYX9+xGK4vb8Bt7fB8D
HPwBVVNP29JcfRM/zYFaSkwkANBJCoY9QMCIt0W9Opm37URba8Q4+g3w5H7y/p9XxGw1sB1O64O5
DHWrn3mulzI23VtYw0WGGMW0KG1FApTxb037xer1MULJjwqtv0rwuIjoUUBQnKCX3fFCD9ZzFods
0fmdSelw896ZqOVgMgio4mF8QLi5L2YSOUebcVK6lpelw+kVIR058XsCYd/1DAJgDT6Wwavf9m+2
HFh2F/b78OybsvYZybZjjpJQzbcsTptoJ+Ycs8qf7jrNnXegy49jSRGNaEgFXCfHBzTMuqlc9tzL
Vrlm/g0zFoSsCVE/yeCLfm3yWjxMQO3NS+HeOA+d6mkBbixvVnsHJJDu5r8jA5k0hu3NW4146v6d
48ydCKAhAKzVWqAFKPAabZ5p5v9wxsJscMO/BD2PRYAgZ/aLr37Lv0fcPzpT9xlaYFcbHANuLThk
Pu/iiy49nxnPXfcg/aNjkmang4ywXkhzIMaxFkNqkzoMeGkYykVGPpPu5R0GvTVPYn1aXazPJU79
kWuzmJrRY3GtbNbMwx0rv/hqueUirbyXFEhm1bKz05+vuspRSc1MahxK2E0XZ7GheNQef/uGL1+F
EsM/v3zr0jX2JhsRu+3liz2GniDh3zYE4v/jgsxzCgneRf/7CB/qmu9AeYPVHOFkm0BrGbMgiMlr
4ogpJFDvBgNW18gzPeKFcHVxuy3++CN/+h2wBhMbJuMM6Jtq7VlFKShheEuyJy6g8g2eiVL8aF09
kmDjdlgYvjvBnOhUjkuRZs9+iebX23hZ4OPkBqhgqAK818QE2LtGGdS5wb5jiP3mOgMSWplAqDEJ
z/BqDB1kwmD7eTD9+/I8hZkh0hKingfrI3IAOh3bNKsYnt4RVKQ6Bq05ykOWUQndMmyzr9WASK3P
LBDhCV3waiTF8E3rScTt+rsUuc9VmQ7/3vCbtR59SjStBUuNzTYMJN3COcfaF2WFhbZnqwEKj6uT
xWi37gLpIH9A7O8L6ruuzVBgHYIWBbM6e/9w4BpJanPEjp2/Zcm7p7Mu+bQeAbGm2Ucwv/okTt0Q
U2CrqmraQYouNbx1bDIUDvMMpOO2QJ++vGziadZJzui4yQf2InJm5ZtcM47LvDAD5/y6YXkF9vl7
Y1MjiKT+6f96AylOLfcUBkJN/X193LI1tDi8xXUcdvEGYidBrB3cg1ilu6ONolcWap67PVMG2hsi
soIvIJ03F23toHNgJM7imi28BQGQWz7U5m0HNMhp4FfANa3X9cDPxAdzhoLfEAlctbsk6DAFS3dh
5PbAJ6pn+Ldu4Tw1epq36GSXJ5f50WiedvObJk9+Dwrw/wGguZxvtW0yBgEMARVU1dn7zbnUj7W3
hOo7gRpAfAdP93AumvtN8nXlFd2t4XJSv/33v9WRYftmLdd4kb/1WRYyivkuXUKoW3v2MUDNFNSg
TuTXiHrqctbOORcV5m8SuZcugmb5JmbhA2QKI1Jzw+FI+w9J+ZxxWUX6gWlIBfNlJLLCgl4t5wxi
eFv/14GO3rYVhAPnO1zlbH5O2yMFlMI79p4hVzB3AaUbd4G/gmbdExslBBs226MMD/p3hLg1KA3p
zXGXCo6FvdF0nswsjo/NTwiTRaM+xLsWZhP7hvl1Rf8r266PergShtYIxZAuSsq0oVelZPcACrHn
I8e0DEYC2iMSjaCeF0u3wVrX73lzJWvvS46tuK0AtiM7qTK/PT2aEY8JT1gJvlFvA+XCff/U+1rU
vtheU8p9KA3V7ZWXyE7CdBApNp1OUixYxT/C7Qvbq2VMfgIxgjRoXaMZ6U43G6d1h1BstnvmT9ej
cZU+K6XZFRE5fFjXp9Y2sBrkGc5WHCCJ1SSIdL+jW2/Qo1ajoYcPKeR6rZHgYNAurWvxugx6dssO
vGHvHnxvZ0aaEzTEJBzuTvvpOc1HUa/Mbgziyf9A9h1qODOU94gmnNOHIxPKQSZlv0pD3BxdHltI
qZ+uGL2fKPw81ViWTAKPHqt7lxZrAyp8V6RKjJXOmi4aIol4grFRC1O1cAPzdVcjOvN26xPIoTBm
6gCkOqa3QR/ZBN9ISuhDO0o/X9W9ZVj4GlqPaSOoYCPCbBzKtaOq+1uuzB+V5+7K92FQ3D88rW8A
AUNsq+kIaR6BWXAOP5t3QEA0IKqijCd9wbOIbKp/pMVIosJsaOO4xU9vqt+51T2tFJN1RydilLjy
or0+2hSf/qFEVRbRR6qdZpms1iZqLJtcBsknz9S8CidAbbeMUI2znH7/pYm/judBu/2+Xv4PoQFy
mI0Igu1UpBzMaIyST+jOJDTqvYm6MzQVHKFJpg0Oqp2hQoBNKpcZo2Zwp9afzdns+BVn+4aoyN9p
vNe/OBeLKeIx8QSTDoEEEfDy2sfdxAMnQKTvLGtH9CCBJXoFUf1gamiQL8WiRYe84pRmXDt/WPM4
uRFdnhsktTmV1MBkG/QnWSaBu8j3Nu2+pJxIouxIB4IT9rSi3iPbH+M5nmHFFC5d0m8tRmjUtl00
HeHgpW3UwE0G0pul6Fyknd4y8bZWoHL+4O6trnImmE4C4g8l2+U4OBwJiMMCPxRLzb5twiP8qNc0
Oa/MY99U9wWJptGh+nHlaNraqxXdFFNyA8ZBnycNdylfoqR78F2yXe9tp5hVKYCvlPEgQjRLNLfb
EmUTd2dsJRhul17iPwnTZgZgPlN8HimlUIC/cGSzgjiIpZFZNySSwTgRZVVHkhQBGVPv2SudrMjC
go5xrSLzpp8VDIr6v0EmZzjEDzx7MbPT+s3qoeJFEMlDVhx8rkGT5xmhbZdaBHZLMSnEeoMp5ly1
ZA3L7kBECSXHHnjIZ067yPOw+IBUF4eo7UnWZcAcFAwJTucwER+PWRr2joSSU8Sv+DEZI6RkFAdv
PV2wGA5BPYl2joEecn0fzks4pJUkIq/XMlHrXw1IT5fBM9ouqE93zkNTCe6caI/bLK72jcrvZJmM
RbfqexSBr3J2Q89djqZns/V8Htg/FP8ieudSNwIiNY//m7Quc9dAm+qSyQ5mKZ8pWKTLz+DT4nah
zxB1gdb2XkYfpQ48+goeLJraZVyrXjZwsqCDp2YUmPJqjtQJmKAiarvv/pty0fpsud2xGJMz07K/
jXPyfwNFVPnbZpeWh5YWpQ20RJWXkBYJDUeVnDCL+NiQIjvoFT5O8y0Xq4SLbypFFoZawuUHoxL5
gUUGCg38WPRNRpL2dOo99eRrHrV3OkYGFrCYOiWy4sU6lZ/uR5vn3/R7hoNarF82JvGLvxPV89Hk
UdzO5gWCAJ5ZZ5uk2y31TTYFpHYafyOJjktQ9lj+5+lFPvUPOyfYuYtILt1MteMCmzdP2En2Bczb
PuI7rvxLnQ1iSsK6i4u03BMQGYxlw+h8KDvgZfZNLEeCwhgYrDcSdVIYeDveGfM/+0hD6qhql9WA
LJ7r5XM4TTEDkRxohYYjLwINn6nCue6LqYisH1FiIw2InAme2aywfne1xj83abcuN9t2XMJ9RcHC
/bV9VfRGV2bM+ZaoRptSmKkiUVfIYHgWeGRlKOBO+iSNBZ0fFzKDVLwdBBKdgg+LYnsnHqoDVCbg
FSjynuro/tpsreYzw3v6ewEqE0REvoC3XJzhbg5NWA8cD9CasId1GPVd+Xw/uyfAx8OLtE7bMTgN
RLVgxN3M8m2yyVndspJXXQJ9awnGIQLrWP+fPdkvBXCTwB63G7STApyxp/0UnN+UYbDz2eRQsHg5
KvjmIwKmr01MTi42HYhk8xDFKzHt/ZSfRCm3oPMxjZAvFEJiqIwWHDyvZSLGxjxz8f9g2/YIVyDE
iAvXaFaBGZDjgZHxk5GQp01/PjOjcnWRgKzPT8N/DarU+0v2moVIN994JOciEl6zxY86blbtl0eF
2Ib99aYZdlIZaoy1zDNhce7jQZL08OApcOc31IVyzb/ol7JyIE/XUeX0Cu0ESYm+5S61uKhITk7b
8YZOB4d426jRaFH5Ht3EohyVh1jy67Mh3Hj/xdwLMeKkF/IfcPMwgjDU9lEotSNQfbUsuE/GIbyI
PDaAXDWJAU/Ao5hCrp9ozgDgf0abnplbbuz94vR1zw7LCsJndX44j4IB4SuOylJUswKnhzPaMOQi
YGitcDw9Zd962fzX2Uc0EhTo6H4AuwxDesQ6BO+q2NZzPezfRNg6WyTU1CETcOu1xZ3SMcX0mNAi
Ic28Ogb6sikdY0681ynzZJrtULXx9JJaCvbdpY7C5Y+/TVBod3yw+Gql/rcQdBqKoUJ7QLtUx+tm
5cPlUqbapxOZXPXUQ+OC8XGjLOBvwpogcOB8QQeWX0GOAYcuRREpRxe6zwB4dNlcslB0479Psvqb
ViDGq+TXO2NZffyW2w1mLxAb2AWk41MjtVJyrsiyxDhhoNqa6cSOK34FU2oum+bidb/1/1cHfIae
IRpM4YWgtXR/nICCsn4fk6TrLfivBnBi3fvF0wG8VlP7yFShBbJ6/KElj0G6jhIHgC5vTb+gFgaM
C2Daou9yhASjPh7n5276QObk38gsaxigTfo4OA0YHgimOQ55QzfqGDd03XyousN+BJvdcoewBn3g
n4Ms22K/gSAGAlcHNHswHVzVCWMLAjE7GmLZQnNSYlFE8r5dNRuMWMrM0PyyyJ1GOqnjBRf6QXBV
Im6+ltaxoP/LqKzWOjo4c4CbiATQp/8Ma9wy1j+PQDnaTBAzv7Hs5c+oZiW52/2NdxymbWHhWCQ6
ijNil0z1fsl/G+/d/ZFRzb9Lems1hD6Xap3VwHTtQKVkG/C415VLVy5Xkrr57uMQ9LgfonGWNuJI
P+in0JGZPX+EnpMJR/iMJ727ywkAunq3H10S1gvYr57/EIfzXjMAFeA0K1sozbEz0U6CvqUon6ko
/1Zgdp5H8r0Phh1jiEjvXdGzFQ/BvI0FB0/cg9iXQZC4IlyRMHKSOLxdf70Aoh8yi0BuQ0Xv5mRQ
5151YMGPNyIjyvDdF4Cb1iGT9yG8v14ThyGiuBFyA8z26c4HlYZhXC6I9XMcjQ+xZwDqnTSqWNfT
/dNsruHD6IEjaochN9VzP1N6uXy6v7CvyjKsrJBa5qaRl4D21fivYC4xtqMncYOaFsDKpO9/7J3p
vRNJVBKFcTiBfRKeomFXZrb5oZHR1W42uzdpJiEgJrHHW9lhMeCL1YlpoBJgHoOrck49G2TOe6jO
3nxE/7A5VGJWz/c/o2JE6ZlPk7YFGUEzcs48LLEsUIj8nYyfbqQrA7YfNXpV4ZCr4tfm/jFrmFB9
C3jfs7qgWsP+kjgJBUEA5YfaZweJ3DoycI0i3lNSsNC/3TkXCerRSVbIHG2YlSUmxExxGd9yplNH
NNYoyqL3aoKVjI6bURG650iSqcAxSqVXi2oj4KeJox0REr2wMgV0xMEkM0biB8EE/uFlLZv1Or7E
c4bOZaeKTa80sGQ8ijndSS6CnPQ13b2QtHhrZfLuej5QSr5ofVrVzsZJhjoI2uBXLtbog9FKoPIc
asA9khOHt9wv48An+1A8LrD5wbBi2qy56Dj32DU9ZkZUnXbTUmkTxQcSJrBdLLRGDOPApoadz24H
qqBuxcgn+Qzz62wHEhc7WDs2tLIElg6QGYLIgEVklZUxrR/OFHmVbLMPUCFPyX2A5z/Zw/xWaaRG
8XUVySGV1gHszAAdfDZz3F2TR6INAinXzTa5LyyLMJWzfskrqsu/8xvbHQFu3SwYgwsrnwIgWYRE
iTIwORQf+BVmOc95HByExLBvo0bDxmDS+mXBSr6zilsCi6eFol28fWs/kCLT6rfVNm3V9seO//ON
FTGljG0a7mbDzVvGwYsiuRy5nJCfD8LnlXkJVzI+yRw8mjR7GcGEUtSseGR/5qW6CqRfR0ulnUK1
24wHrW7dAJpuoiaJzQpPl0xSv3zQROg0doR6xRv/92faSN3leLAV+xN2VCOhLbVUzXCWxT0oIHev
RLJkuT4Ei+XWiLZe/EbRXhnpWR47WxPBJpsL40cn/pOS5MzXD2s4+LqVQvhlDGaQCj3JTvBU+qh/
CTlDk7uMl3oSoCuKqWM2RgLnI0dSWZ3vUDhh/i4XhrNNxCrP12cI4qxD2PLEKlbs3ve9jMIMyMGq
ogqPn6QfjBYZinlUbOxuOlRKztDTyTGYthIumVRT6rdqC19wN+Ov+vm4c4564i9jaA2nahdxECuQ
Txy722uZyUtQCMUoj5GpGlAZNZ8oArlmJRj4uWoPlz379xbQUecw5CrvG7fZYtpxnhxA3bUm0jPm
uEt3CjuCGhdoCIsYpe7ycmv/Vy0WgbwZ8SvTv4a2pt5jsllIuMOMt9GB7N8Xokdv+KnkHzU3yQhN
JXWJXauCueV6hHtL7NUj+XXGQ4NY7edkDlPLggtSUdZccO6MOiV4XbQVot5PLH4FEqS0rQzhvJ5J
3IRBUUr0Oef4QJc2CirMRoC0goULa6oF5x6I4AUSPokqGsrzRAlYMVTmFntT7tgOkrVzBrm4urA7
QV1jW3KBBRKu3iTzsJmEu2TeNiDcDviALBDuvP56Z89wUtE/inWNEkvkJaqyIMSI3iP+KXTS+xrG
rZ/N7LOtYgkuu6E8YVRuiFw34V/i06EKELdlH3aq4Far2I/Pjk2b37MVJFhIRMtF0EZKb+4Wcm1S
08e8H/6lPZB4TacAu1YqrVtCb2IJ/0xCvir3DCT5LfsO4KqYz17LnQi5NbwXBgMwbVpmQu8T8s+M
akhBMLxNLnxQh5kG6FMBoHDeBPJmmXFT7OjkTj0PwfKTrWHWJFX4rOgvF3IGi0e4k7iY07glGB5W
ZEl/n2CYzM8YGsy+JRP4Tc0lN9sC5U+qsEN746MnUJ4bXzpl+FBGB7jgSAmUTwcVGnSKnt7aaKCO
w1BUW2YOXLXv2ChKZkehG8y5uCFWXtI6+QhTOX5HURSEndOAWgFqzkZ/HIEWkUB+x+Lk+ql5Rn/7
tTw6/14FNdv4ZgXMK8lJaXuDZS6/HQDn7GuRc7fkiw9UmX7a8WxOdiIItw3mE6HgEj2Dii9TWQG5
XkwE6nQ9j4O0AR7w8cIG74wNBvXUOAUTVZDs5u7AYzcZUMRzQz276PowgP30l1RUHrMtnBJ3jjBL
YoaNU+C0wUoDfiSYaIrhdKgkEvly53iR+iOFGHqPLcRDVv3xFqvn14iBXD+Xz60WHpeSTH2+9Z6z
VBV5beXUdQK9jrAa4tUCWuFNe8ELnLFy3dN0lwGHfUx60EzEdXYT+oG77l77cLOsKnMUZLy4E49Q
Wk6Ilyx+jjk9+phV9c+3CwdVCifc/XqDKnw3QxbHJ5mJ0yY6y8y7c2k+hj9pXYSxlwMSeDWSw7nx
VCQIHZ+c3KNlPvginlQ0yrnMou8mYb66SLKKttHgYPTVE4G4WwnQBTr7U5HniNuKnhvHtZ0cfeUv
RR6zXMvW6ffLBYU0t16C16rgn3gK38e38gxuVpFuk9hNLKdpkqJGUfKU2Sec5YGktq2rnZPEfEqM
+Le7nBhnhEpLHWQuBAJQB9pf9i6ZokwktsslhWBcRMxxcpIDohlRtN7Chva9H5NuxNWUZdRFj2ny
Wt4Y/Txiw7fST4ZJrcw2TF1p8n+I9wfpWlAHc4tMrDyqEBVLMKX63HVhJNe9YEivoRKZLdG6WCG4
Q7gn3GRL3bPgCMABW9VYeFi85znpGXZEwqm0Ogtcm0LFw7sBe8hmmOsQB9ADg6AZhEUcmRW7RdcP
HTPTUx3jFP99Xwzc/04nLKGJ8Fwc4QuJjx0yci/Q4vZ3pHpaEQkzqBKVKXL+NdVl5PiSaIE9JDAz
VVdst8m2ZAKcj2Qx+u2rYalDvJRHpnrFZnit0Bq9PTUjD1Eq7laxzRi7mzoDEPt76kyCVcrupGWW
i6L+pHMdtj7rU6bQjJjI+w3VTd56TURTzgX4iZV8j+AZkHTCjDKZV8Hg1ObwxAX0unzo9T4zybcJ
m8cOvfyczpN2HZbqQ3AduI63eIi2viCYC7hOr6WbzCumK9PkwO7IQntHdSomuukbstmTPSdoG6Ph
oFWnkTEbmJ8SN4U/Yk45pIhPdTp/7TanNzCrHo0mgyPBmTQBK7eKXHR6gcXGGpFmJfJqvzbBX+az
OWflZh2PUPdcKCzi28HVJt+RC4LMPkBgTEXqvOEA5pcvMuiTbRXE/uYsnsGiYoJeisk2cEN/4OZm
4UePdPpZJrekImuk7XjDmq2v6MVQl7vh5f25WCOlRttm7aY7lanA3s+VxhYGx4aFKsbcD48V6BW2
V1A1ZmvKLHWil0/OpY65WMR+Md/wkVJkxQCFWT6wVYZp4JJ5tDbetAFAOQ9Y1g2m6IxvivKcdy8S
l4Oc4s5VzlQ4cQ8R32fAUmH7NeXV9hWlLZGhPr3plYW/73J1mA00VUGF7vcR0cstTGxhs+J4LpC2
dngGx+/X5JDZ2XNJUbXiBR7v1J8Lyl0iBg7g15GRhxmjrpCcbsqF+5BYMeeExMJvcxdeILiJN1Yq
BewQUO7PUhdB0fN0hnw6MTdcQxqt1uAim+gQfFdZTi8c9bncW9YdP8zaWbKGhs/Ka7NaDFSiDEz2
zlZUkmVLsGUFQ41T3x7jquqoS8nQPtu1Y1POI0rwLNAZVANzTLyYF6HKBrc699cSBHCRWhWFA/x3
znqf7qwAP2TZA5Z7gThClq5Jr1uKDKp1FaQNp4T53gShrF5HlAz0Ge3WVx46rstXXT5Hj6sRQq2o
onwpbQ5VYSlGh2rEPfdqZ41/NLwUpolNecXPXrBKyaRs/EGORrbu+ZLMp9Wk9CMOWLTUPP8/O94s
54QP2Hoq5Ikr7eDYOj34XjWP4OQZZghPY4Y5mDQjjatpL7pVkRDdMsaZvNi8QqMZlRUIY4sRnhuc
nUVN6hFov7ucJbit+VoBvE8f+qA10vE0J554RXHCf4VjmhBKOVTAdBAf/TtJlb1TtxBQrV5225fT
og7/JupGfGZEvvSi+f5km54y4479LGHi9BkP4pEgCTADPUP6n6rcwNcNiUm0jcMMg+t2lPxx66lu
gSLTKKPmZo7b7MdBjUOowcFHB7j+KBOOF3EQLvGjNoRxEswweSOWj0F0sVBQBoCb0z1EVFyb3JkL
rpi7Hjhtxxuwd1jhLToCNioSMmEXtXL6WiiciSVBie3dc0oRz0gK46TocsYx+Slahm0IP46mRQzK
jms+CcBJ9ex+18t9D6arWuwj/ftRP/+oNGec1J4xBue8wS+jTm6y2eI7D+9xLX8tmwtm3owe5oXd
KZSLCCoTWT66vTmJGi+GzFh8t0TXewS5MAkJsH0287DQ/khw+NJJRa9Cwg0mbuWz2VKU2ipSQl3P
RpnriZp6J9Fwg7NMzoPzXqY3cHSkTEfw+TQ7nRJWTZLwE2BotWqCpK3cZQX2BMOsohDlQihlw5Qd
Jb2NtkXIX1AVeGyJ9W4Vix40Q+Goy5uw90X2OPyEKX9qOJG1I8O5f+2ehRoaFpqY1N3m9ogy50eU
KAZUDNrOP9MSIk9VAcPQcq0Nrfix2gkvuJYuYwOEJ3NDtFlktF937IKWl3+aIHIKsr1z1jNqH6jj
/jdF605vCwhV9Nmp6fzLoVmyquKA4mJ1dyDnVR5N8gPJwdi472Hy5U20SkdVtXlyBdHDiN0aDsbI
SwFnMMjysVMMf8n/+9No09fRL1duMIMo9j3zo0CVOtfix44dNTLrwspAzzxORVWITgE6+WUakuVU
17Db0Gd485eqnrTkmeaystlPzX30uTuEt+ZBxiY6wvXo+LPRsL2oq5MYnfpV/jnWUA6cBchwAa2d
YWYMOKexgwxcMkxtXIFw5wfiyjlG9Ohf2ujHczPIbIPtxRj0GOHqYukhNXhvwCH5TArIE2kORH3d
50u8Ze3if0S3HYrPETtui4yQs214PMrFrtAAj0ngBoK/wmYjB9BOpTIt9o6NT6Ok/tG9Tb3rHZKh
sL5jaV6EgyVSJPwOS4UvqK+f4j9t2N3xJYu5N1b6m1SdSBHfT+qEDuDlO+SfOfsIKkBq1kBGFYj2
xgxiI/Q+4q+EE06TxTPfeF3LTTcKT7/kp5YDCSqpdQdD2Fg+zpyRYIJ7CrIlFW3vOmeTxJOA7Y8l
/OT2OX4bosllpfbOo9AkW7yix26ocOglyM1qeShbY28t5itXn3aiwNtj6do/c/3i1ZyTi7mFtjrf
zfmeB71n+pHYnW99haKxjZInS1xz9lY6/yFak9G08xy3lTTr9w/6TDphgjk5xNiGkFiXFjZ+mGCu
EHuiHTyiM1zh/7d1lOZOvuVmcEL5j0ZpK7OG91Nhe73CFaYvV4Od1k2O2ToBr91ynJ3qh1VWFoN4
jv0WzWSon+Rjyu61HvZxofZm/F1OaqqeZcp+t3oU2+CTP8kaL5/h10fmJeZsXdnZjqxnIF7E9U0+
lyJwz2exb0E9YxeAXA1R5KwWd0H5kikHRTUkG2nPhSMRWf8trUd6YhHrJ9jbgZU5khN6CsfDGF6E
V8jPoRtdNLMiFqPGm+RdYS3ROAHwffkYkudiNPDoPVgtnKz5PnZUJkDtgWupVAS4XWRedDSxRBb5
0fUAjLBDN6WDPZG6hVMbHy/ZryOn5VvxtDKL/nxYaYqN2muhxXtFDPUkSIhAVmV3NNBQeXowm6OI
BKXGw0lEaqEQ8lKDc5hHhF5RUliTs+bGhlOCu5Yf9yxnpgTv0PtFPe8tYOheJZftxZdJ7pyZ+E3s
itC3TS/uwqM804xRb7o0fjTnEkdMU9CwDjl0h//T2I8qpkhp1H86Cye0WEQh9kbQ1ilvqejFt0IM
nguBSgGGrNHAsIIvEkgNQWUDAQP0Tqyxx0Ucy5/6TEDm3iTpQJdIqpO65CuH8MBGPK9D7oud1rKE
DqUfxtMHV4U/GIdWHicDqJpvGpotjppKaTstE7He7hVR9t+E5z+k/PsXu+G3hSj0leTE2a3tr5En
Td4avxQHvGX2ZSWf0pabBIUPPtIN8lC5nEMzarGVW5a/ZkSCSeb23Zt2lBY0EqTvnie28ZAfUUnd
rmKAJJjz3FiDg3i1ZwRvQF1gsUyuw2bC1s4ZDC6l1BV0C2IEK6NpBLDenQiUVehSZjF5zJOqVJVc
ZTpQfcFcDvcGp8J+ZJrDkiqAWrJu1RElSTb4vSO9EgKrulp/hQoGZ04NPYE4HucUPCvCpApI4TwZ
6cZ9tEC1cIXxWEPgMQG5odpbahZk0/5hMtKJvXvrBm6m8Qn4cjC9uMY9XPtMMLmRTTeGtcNDthnQ
+D35gzsvRtIs6tu4We+T5U7++8TBjRkW1EG7SPKhrx2XNjfodXzcnYvGLaU3fvsITETPzWuXwBB1
EUc2Y4DNazVqsF9UHW16ZGtHxfjIyxQCLbAo4B8hD43CZBcg/1+1VspAFaRwK8mY4v37gs7WAnS5
Gecw9jX6TYvtPnMzZhuUEQG7+W3um7IQGrL8N+dIwnd9qq6bDVzDMhpdr3M3XUfJrCroDbyMshjq
capwe8UvAcPyYsMaKWuXeFkWbYFvD7BDqJUvgYUnmT5OL/UEDT3hFoyUvMyQKfs4GzAvMBXfmq2/
3mLTcAMIlzFRBSdV6xel/mrMsiOCbckmTz3sBOBxbSp7/cVQLGlxzilTezcNgUQkS6Ut+r+4Jba3
eRjfl+oYke2qRkCsM3vZbgLcoBqp/lo/Bnb/y0arkmQNXYF8//EyYWD02E4tTh1WLq30y6eKhpip
hoC+gbLfepYF9TE/es8oYGe2xIHp2p1MXFkJG5VtcA0gXA+wJD0v8RzIHw4ybA8uR+/mk3gMR0DL
zqz6VszB50XbQPwcl8ksHHYr4h2fXHaelr8Xj9y8pHzgMi0q+wddWKY5gBCyedYto89UDnStnSOL
iPWt60Fk1PZR1pAia/U8mLPIhsI9TdJSe57w1X7Ra+7JmEgLyHk8Be5EX0FXdQ8ZcSf+VkfEgvNH
RMpJf3mF9VvXm6Fnq5xcshjau6tCywdcT7EQU1njU0/ueBlVZE4twaJeMGEYXEflvE/yCcQkyfMz
QELIwNMYpLiigGRmfDYsSYcXwbIFG9MiXmL/DfTpnOE40eBhzK6kYKJTKz2wsNbewxKiRdwR+k8T
9nEgMUJr8Q+SW7AQMs667q8gEEoLzXoU6Iuyr78dkfv40/BV1HeEC6aPNURyrPunRCybE5Gcc7/K
oL39NGJl4y2dfsgGuEPji/dGzm+hwI4p2dtZSo/MEOjUMS00UuK9MB1q4XCrXUQxL5PNwGFkVIWr
pR4kUu5neTAzp7iyJ8dNr7LZOWmjsjnXVs8XQDBP55eGnkHtKnKskdKsNQVZDu2WqvSvEdQLQjLM
9Q0VepUAUg9oSyQunq+i7bt9skkHaDZ4Ft1jrrHDS8YaAXaZEMtpoWnNLASfGWiKxTDtVH+TqW15
CWSB++oKPWXAtPXFhg5yMcPI8pCnP1NPmU/jpM2LGEaV0WjY0OoL8FFV0zKXowKJ4OzkYNzl5M2A
1IoF5YRyoKcbro6tLhNcGpDiAMGXmkyjG+JeqE42ZwwaozayIi3RIcqr+efgwJXSmb6ps3UDdXgH
+093IoWASj45zx71HVFRM7cbwdAogWfBGr8QveHyL8zoKx1zIP9eXjg5Yn/TG2xyTnr+SFsWwopJ
qOTt0CxBcpmFKpu70ME2axbj2ItFcUxKkyfzxAKejHUeWjnR9qb7dTX45hVjtloUUsdLaWABbxAU
Dgq8ZouT5z9Xnz/+g/V2rrDeo1pDmlFmtNVTMoWpN7l6WtzHPEBGZqSA0qZQOwuLfCe0NxCmYWVD
hFAigOnnWqPkB74rQsNAa9yuxll2jkxJD6zFUhZ4oY9jhop7yVkzMBYq1XmXUOluWz/cuITM6m4T
bXaE9iHoOcCIdCOgDODCEGoZTSPzqDuQZO5a4GvUQaV38W8zunMZfpX3x/Suc4GK0458JpiK9l6R
B5CbxzKTGRAofg0l1Trn0ix/fTBBVre4wu+zSuTso92JiqgLP/exaWqvCnFakkksdi3nJD2IIWEm
8TmDPNCFEHTED39xAx0B0q76bGpd/S7AaB/8L6Y5BvpQxlx1Ek4hrgHJu54r+vWWXljlfwgL9VXg
OwmlPLGGtZKuEn5/DxNot0SDoXAp5cSNMH6N83FNdS4A4wJa5DCpndX0XsvHQT1eDwqGhaQ5RK9a
15H1SLHDDg5e3z4GJX2MZrB9gfwD3OZFsac7O6uJNmnCJg7TJl9UYAX7jG16Z1sXwTTp2JDM4rnj
IgHgx4YlTzQkknbXp1iwGTuUd1wfj86qdh+zQrl3zGPZqpsUkhu/MP/MAuIsKpG/baktalaH7aFs
lH3TIQW2WPvxuXL+992mq50MyAFtd54Q0EAEAEC7nWn4K54t1wI8DKOi1Brzfgnrz43wjeHYPdbM
NloLY/T3jesZcSA0zPyj782oZYFoF454v2btOslnaELAGNvoqAPw8/g5s9cLtoKnIO6o7nZGfuIP
/apbjtgHROEB3N7MNr86ObLLysjTqMf6yB39EhM+cga2rB0HjFjD0NxKMfOi31Hb3qhMF9KaaYar
JqKDucjBW9kqwkt7HI4CttNFPpS8Ii9yPkGovd1h2iOIVesi6S8px/GJXoQdhzqjKwm+Wg+ckRdE
xnWTt2+oOmy0TX9/9EvBT6msjGsDweL7gOJQUymMgPQy6vrh6uyy/97UNny/XQO414ysP2epYAzL
3NxyVhPpkCTtF0uM8KwdDJJ2zBkGc4W7UDPfzYfw1FFHPKFIwUk0v/25nVcZZk/VXFcqaYv59u4f
JTZ0QzA9XSqfDUjtdtEEJMB3Ua1dP4sThlUN/32y9u/+ygShjKyOiaJH1i1km2Hn2fmikv1ye0Nn
UzHSFLkt/fcHLUXy2fsKIDEsN7DModU5X2F95heald4NovbWxjPDcC6heH65W8qDOBWFklI8xyfg
rLdKsbuYuHuUITItmDcPyFtQsGhs2M3mklc7kRuvLO8fbUUE6oS2LYBRiXDrc1oTABsCSBuyNJbQ
euNc62eerrViyL/2IDATM+YWkTfGx6foumaiQASmM/m0YO3CXoII7Sd8TVP1bW3sBi9mJGpNRzkw
Q2QBDBHkKP+V7Ga7/gGI6RavbgMpYMz1s3v34+eWo+uOUDksLOkozLP4moFvcuurV2+OzlXNKaEK
GpjKLJ7MAXpR083xgshUcB+FlK0XLy5fAoEXqH0upbRtpqRXPxT30B0JWbmwGvOcNbLHHRHnLR4n
IxptOYYrT8wi+8nz+7HKfbKwOLpBZQeqRauTc4gQBs9oDVIsPpXppfvMrYIjpazAoekrqJ2lUAe6
JbQIZLNCh0JjmRiX5UN8meMwXPkJtMSdNrB20iAwNxAsTEDoZz2MQTznTKS4IBoVbbb8oD62rC5/
1Lls4RgK+BE58BFEigqStEd1W67TmjUoKsnA7Rv40nEsjRff+7QDcbTAWRSLhzWFwpeEG2DsC3Y2
4TsQgU8YMBNdCexbzQO0IJW/YtOHoG1mcROsdD3iemxLXdYmxXF1yLhNC3V8v3vpFnQXiXYuUf6w
VO9xB7r/7+22mJgbaGX8VSeZo8OWOwjAlKeBrYvNV3zb8m8Qzl7mXABThiNAJwP5rnnyt6yzJefZ
JZsQZP+4JGo3g2jj1hvBQxnj3+LeGzA2uGfarsnnWK7Sul3D9beAFIaaZ9JjOzcAIlp6jOJ8jKZN
aaGPAIYE1/dw8y8RDyrYYDObgMvEifFeeTfCkngkw8SpamhYJtJrpTWRuQkg/VeQTqSlC5hc/5K/
VauRuJbe4In10YWo85S/ly7L3IbSx1LLvHbZBzAtk67qlS17EVPjTa3W36wI9gFO3Lr2qH3G5EZ4
ekPXrYX5eXXOLmDIA93k3qfb1+uzBdzB0/Dop0gwNBXeaIPFg/Cb0/mdfL7PX1lVqxkkBHZTiDej
LPbN6sh62JcrqY3O+txQMRyETXQkp2BSy3a8ppTWdMsj8hyyaEyz4bo0TyBEm8AEGERReC7l2stz
FoqkwtwRGZpM+/CoSJQMYL9gCovRPp8FNOyETzNDmTnmlBcMqfBtqn8MCoLm451qoix4edpn/yur
WuQj9g4kbDxZXD006nO43kdGkXqX9K3bSQkJc1IGPnCDQkSM76C3e38grzacVZVnJgOQCPrBJGFY
Tvrbl6zTtVLrbPm+62PQ7fQ3CuTy0Is8EvARv5FAiZZCxx3RzEkK6EEAMdfZ9nCl+2Xyb/NtNegQ
lFWNmSm8qxH6LZgIsDxbSwhE6kNd8g3axgwZog3+/FCC83VrFv8lCFIdo5iw1YgPv0SJA12Bsi/b
59+CvP1YaNyO/YXK5h42kuaVhNqggBPzs7dyxcVDSDathtLxT/xExaNGRUxRSdK7e6CK8IgTbgOw
Fp1mxjhhfwZKMpqDLRXKCAUpFbadYbIv4YDtqpbhLXYj8Jt9wAvPqXxA3vT7hCg+rSP+QIxdE4wv
G84HhKlkWiO3XNwM46qFNQHUKdzrYQvwwU+tJ5iScP7m65oyBsivwfJQXEJjUiAOF7KcAKYcQRrj
JalT1UY+XKPLJlwHoCrR/c6WU0xYofPoFta3z7HTEhU8u5UPIOmhJZ9KBQ8LvPYoqaD41nhYV7W8
UsGd4iM6gkCAGS/A9h2OexctFV6K1/H23MEAyXR0PqL/TYW3cu3qsxXO8BW0JP+hm+Pmz/LtO69i
lziXVJZ+3Cp8tSKp+oHF9Y2+8CROiwnvUBCmez48lb2ygsEF3xrMpAOSyraiy7lt9+VRABgk3lsA
Xr3X8LaWI/oG894S89q+ShVGtnu5CCLr411EUKihuWVCVsK6liHVaZFZUpYRp6xG3gPv9GSy6xGP
53N9r0yfsHJBDBL2O49PpiQZuIIarOAFVZ70bHs51D17oam2FRe/KmtvxnWBKRFHgXRdg7PjZEKI
3RmP0YmR2cRWeIV7EjybkZUTyZePSId4KMGXeDpT8axbt1ovNw2aGPx1X2kOXHss34vcBID78W5c
YK2Utz6KahyL6GO6aNOZvtMPnl5+n5bLeQBDZQYQwNrGL1bVj2vn8ht7nNEqzskbW5j5PP2EGMeR
3fOXfhDKCd01nxn2fUMBNEOsJKgpFZMFeVhBqSosXw+vFzOBzCTwoVeEgmXx99kVKZ4ate3Jvftf
XZu2rMVsF3zWhST45Ozv4IWSw47eBfbLRORpSulTIwfSx/G0WXEaw/37vkXLCp6UUzqMCUibM67Q
mkpj/Mm3SYn5hudQ3mG4R0QW/IY2GntejK0A/3MOmC5q1gT3kdMAUjPZeHxxuRuYwdwxa93gd41r
srNEecNZVKqoTwa6YXwk6wafBA2iwNr80BXgEq0SlFS113Uuchlv5JVn1Y0IKJ7Tt0f/xR/IWwZO
Cttgg0/uVEq6/E+rMkzFB4jFGLireb8gwgm9B4pLjybay9k1cONVXivXDJpJTSC9FCP5WVCFeMqM
gvkJyxVBRX8SmUSrxY8ynXOHslDxVKDSb7kA/GS1qNwAzs1pSutcL0/z0OeRRjFM3uNuU31fqhqn
hL9OnB3DMuSWIVbOznD9bRet+fkgzivimd0EUzVrkoswY5R1WAdyWh57fAc4lX4cVNYfQjvMaXnz
LF8CYluo2Rh0MLJKE8C7vCZd6MBOS1I1USp2GvEZGoZ4g0ChlF+PitX3hv1PuR4Ypx3PPIJSqvwR
d6BgHJxWC3L3igehCXcMSrLRdpjoO+kcLcu4Cqmmqb6dIWhXY/0kMCgplEvHCF8p8J8/J4loqJhi
SQGafH2Xs43PvQiiF57FrvV5WrRzbBZZQqZhcJ8yuTIvl8Fc61sP98qy6YjEK9DYX4JHfvAhRczA
hxa9g/7I4xkq/H7EepIsSh/Hw4FNuLSOa8XKHSe0TEizLB1rAx7fnWKLa7ZU0Lf8GyqsvYKGN/D2
JcnyO37gaCfedZNVJlviI6zrcXk5073bHJYvNXgBuT7I+x43gH+02ZVE9mbX2hy3yUTbe6T3yLxv
bPWT5E5t17DmSREp/Vjnxniw+784sY/ZUkZz0pqObTh7JR9a96oNBhS4DzhRnXb5CceETwElEgBk
y6GDTaClDpYrSFWMEdPT6AA1GbIbu9QzCzKX4829+IM0zug9G4tYfJIrOMih1T7ZscoHMqdRv7DP
l6S9Cu/MnKpCAImzDXZzD4leYdnGxhi4NGR52VslwcbHhLEjbuqIlVZiFchL3d7ds6er8hJyD2V4
s8QWhGEiB7dkeOl3TbOiFrVZmVSLB5DXcAf2P7/afeLnxC6c6FTpib+SS+g2F7ozvG2xRoiGHz/1
DK8gr32Tis9HWOL9fB/vHrBSRCVTg2pZ+hzJ1UWXZlfbFaLMWsu/9+iL7EYAJQEK/ZcL2L19LmLM
c+AHZHXlZPt0PePzehspWU3hQQ2jnUjJUveSW7uZVGjG/zjoAZgpy13522EWD0wOAbHcnJU3Ai2r
zSbIJV3mwcrmwaLGsYmLYXfxdO9/59zISl1IkVFwHJpdNPaeDEegUGdpno1gq6OIYLg/Y1I8D6p5
0pF/Zgeo/VjyXfTkGAj7aukyZNcaiWOkH3fbKYFiPhQyxOgK9GbSnX2FsOq54k59A6yF8mwwFhMX
rpbQFEbFxtdDkaFwr/38Zic79ZnS1q5PBfv1m6JCYWfpTfo8DkP/YJ4KuPHxxrM9FAQBLYhN93Jl
3M+c0N4UsyPCsPTfwf3DRTAtPXb9VHrsGt0DqT/Y2PvgWDuxKuxE/qOgPi5W4GJ3kb5YHpbJfIK5
7X/VMW4GZlVXtILhEpAN+YxnJIEFjlC9ocwaW2lst6ATM+z2DTVhAnAHS5BXjokBzbsyx8ux3LM8
vawVIAUl8MBRsdkcAQY9KGp39VEH4wSHnT0vXPUdVBdGbMCi1Fnl4lDc9hZi7pMyk6ZnjktO67oh
wWOWLDO6vnOLAtyLIzId6kA7RjILUqXJOKAi4zWdRmfFh8InnUlBkSwlXIlJsO7q42uQUn7vn0WJ
6+jo+8Iwzqcu4aJ5dQ6OKOjkCUxEC4M7eW27VTFFLTVniS4WPJ8MlY0wezpmBku/0GP6CxTLU/QV
m3ZAeloy4z/Ia9TubRe7n7+c4woDgLYIti2fQjhztpPFti3aBj9Yb9ZNQfyl6FnaMxVZLjbtWEPx
D1KFqyBy9diKxSjLH+byUsw/z9aw990pDpWNrtIf2mcWad9bjoa/glP8OJq+lk2YHBW5kDhLreWX
tZNiIqWn0OUlzgf3idMpgVLinlL+L8xTDji8Qry/IK6tpmtv+Hc+f2UOGeWYqwjf0U6tymcridOi
DMdxmMiIjj+SARDuy8sGyB4EF8AIuoYgXCngfqGziPBlNPzYnbxhMrAPNJHsPnTHuvthIY4OQDAU
g0yYgkCEZylTlJoalG5WgGn5n4UZaYIsWC6RnPQrX/IFf/HK38vEGMwZFltcxX+Rfh62OyWjdOjT
Z/7eEy6mmyoGcmK8gaTYLOFOV1yJMu+O6nIbNl59Gtkki/XN4jGCf3Q+JUe3fPUN7WtJ7mzxGYU+
A6uL5mePG+H5MlfKY4hdNl0OG1pGph1qwKsfm1+y3FY2YZ9Vo7Qwt1fT3CblO19ZHmVAm2Z1E/Vg
7/sZnV6aDRqYkDFzkp5C6CWmxJsT2qnufszzlps/xgwL4JS0F3JFPxd7iZaBfcOs8S/q2CP6DVLw
Jz3ybSWq+cB2xxXQvgf6VqBxoX0umyZG3JpdFujtoGickHeOh4SGTFIoSYRm6Ww3i5a6Rkv2fwZr
/fAxqx314NvqgcleUOky9VSSYiCNBvPN+oYxDKYM3bUwe4RfZcnN5PZHlBLKdof13hLptsUqQMd+
xlckQOpNmIEZSwENZt4gmBcWzr4Pikp7J935Jz1AlSRoC41g3PDz29q5I5ENA1Zt+DzrZ1wbpJtG
4x+RpZYJjRw0U2NCPDIzWHmwWiBJLJ41Qtyz+ClkEeSTqRsxow5wrYBcWvrY6Af1ENeoJZ/NDQAH
KdrR46DfHeYPwcgAFLj7i8J27ZvT+t8PEWzvTqrTiE6Jp4DRU9/guLzG/m2P2tqZTMP4015Bg36e
7xTgbRUrAAnlaB4USlQB1rvmTbpQiCK5CumHOqnibBk3N9oofedlGmndBTvCe7jneg9jiF3g4QjD
gT6fN3unSdUPhkUsm/EQiBp0Y8VMB2hU1ibwsIKBK7eRzoAWnYutM9HkyWHuHIZLReyA2XTxJv1T
7o72ryJC8Pg+pOPy35iVNyeHlu+HXreTiqC+nK871NT9msS5OGl4o9lhdGmIB1vS/oe1JzAwZ4Zf
jQ4NZ8pY9+zJ3/EYnp8/XCrhAApmTHNyo/4KsunxF0aY2F04kNTpFoM96d6fcUGEiyRsN8wRHXZt
xz4kXDqkXcESNCSp0VHQrpXOSMmmfORZopbV3JN0/fDmhPQJ6PhN8Sp/Bo2OA5eoSLSLQHmCgUxQ
7K1C86R5YFhFt7uJ6Vj00KwtonCAaIScl3epfLYkl3igsOMJRQpfiVG70hA7wYrsxLH6AKdE36aN
Rvah0H9HrCCr3H+rYS1tgQzXTjQgH9tUDAzV8B5b2BuaZbpRxpBUASYAtWPATWhhko1MO58PA2Bz
KdKlacm/iL9IH0fnPm+pqaqz5fE4BKxdwX4cml6TmgjFZDQebKjlXf3nrgGKYMMXyYfdGSB4dN+3
9fNuU/2F5FjCBOrK0zR53BD46NqmFSyK952xRL/+vQqXOwubI4LHF+dE1y7sZzxTnT+f2f5fGi9v
A2dHOvva9XeXTfQ0AQycFRE01ZWSpjicrCtQ7HjfSDlNS3xoSCRuSUU2NxG7SH+9+8vQTkOcgEbP
H+gTRMDX3myIlkgJDqv2ozHPzua2z2VYpoGF/Q94DAt37eFOueake48VU/4+jroTZgC3NPtzgx/h
AFhH9CTNIUoxyDSXyYrgDym9VM0BsY0GYQ1QcbJpDBnk7xgFepTjGojzwFijpUHqcAYihDB/DnU5
+BAc7CYZJpN1r/T5E121F1khtTcuLrB/cSmKUIV40Hs4bYPPQZEAA7oi2KTEZd5R7w2qDIMRgzqL
s1jjmXp3BbWDMX/Yxx5u7/CwcCzMwXSw6i05oxXhYph6rPApNClhRNHaO5QTeu+1XKPS/egO/CRF
y/nR/C5Y+vREI2FNZB1P628cjrZNddfhuB3XdleGTmPYwImby2DgAUYvjxathhHz3eHd3+PXHWwI
W0yziCZ5EvCm37mxxrs5CpqfSSiQgGM8xKLiV9PCaVZqQQNY0+7j42QoJegd6/H+83i8/X9PPOGh
iBCVS6SjpzrXSCvpysG49BFebr9TCkzGTfyU9ZBkGL/xiVT2EYoXazzmoGJiCv41mxUBO6alruvN
aC6ztLrfzRuOludSIB+XmdBlQpFP36a6p3gOakuziptF20jqSKxmC3La59B8Qz0dc41FIlsgGP/U
/jErk99czOGIer+CY4/G5qujiE08/cqQr309GZDzcPvcXGf1nqFOxgJFgs04DB/6whvl8ATrK889
85oITiEzNigl8cEG3vXZxvr5GpKoNhElAd6UCvOYt87xnEVJK0VuXfc63gRLIYD1I+xgzSEUDJka
8OHMaauiYyo+dlTiZf9s4CjEDhaxW8WuHWEtgRh6NkzkQwX+VqJcKxXAIWlDkJRd4U+Q0ZQvU/qJ
kONMFDGXjpmDEFGe6qJIJWFXuP44F32q4X18CHsOYhDIcjcmdAXnqrd8wyvp3wnM1Q0A+bMyEbDp
LqumR2HjBRm6d819QE4arjzmfZPUk6ohAz7bAYHJzrmadZZr7+Wxh3b4Ffl7NQ9fZjD5UXmuKNIu
X7mvaIlknD7RIO1m6NnRhAs0HF0nH4u5rQ3aOvvZmpCuOxrNczeh52m6sTnvuSCepJTPPJRaBqku
I+VZsTE5XOA826BKQvJ+mO3hf9C/QPf/SnnWU/6hIQIRUEecmw6Z6bgw7TZTwXNo0WbTdkU1Qc1P
Q0xBzNnWSbcGv15m2CuL1d8xbONd6/XuFF3zCfeGanLrkRRNCsXQNq0mJsZN2qOTBEU1BzYQNR0f
3Mkra04mfz/LdqRrmupR6YpZr+CILNaEVncRnqC1D4mrKESoxN0Z26JPRZIru8vBy4ANrAIkZgS5
FEaOadRtYIY7utRa44RJosJrZz7cqKX2jWQ+dzwVUi238KWwUxA8BIjxsrjcx9R26kkWIcix/HUb
t8kNNetyfXx3ZInfAxZ0qBVF9IWAXCHl3xJyofvsGum8fjrlSNfhv+tXYuxpoaTd/k6q5DFtktEN
4FRz1M49lhRPECLlAh9IttYZfbgfN5NyDFKY+cepgj2or8dccIZdqpqScXFNlwynpO3S1JVOrNjC
UnZr3b1aWHhQFuVf6qvdsCwFbNifEZeAw6pP9+RqUDpC1lhNs1fuiplmQCAb7haCeQPZtmyiK0jJ
8taDTN3zVIJ/TUSfdNGxDMBN+33M99xN2MnhubnPiHjXNg9o/35KmQlnKLJCEQIseTkqgiaffT/1
byhIWCfyR6VBa8VqRQ1U/hR90Xst5FiiwKhAe0M8tatH7iuUtL9zLdlmxvZt37bquSc++P+euFMN
QlDMFPfiQ8/7/BXLUxWOTRJAu8nYjVImKilYGz7VcSqrrRaRcbzuK8CXlhm+4MwK2q8cKh//I3dn
KyhkRcmb9/tGvW1+9CVCJw+Zz6MMyT6tBBk6HixRem+3JP+nvECbDBMRtb7fCcEsXkcB74Vipl4u
hTHB3+xK0MMVinHQ4Un+N7igvW54VEOvdLa1K0uJ90SnvUeRsiB6rFUEsCEQPZ8RG9wwT6/YHpFu
bDjUgbOPrU0U/QMv9GF940JGiRDbeU8LKVyPy9sob6usadHtkffJoBu0p/62ltdunYNCeOjqL36O
oX5xtFqyVQKjnQJwlJeFzpy1MigTUd7Q7pxXdwINHhQQLsntzvJLR8NpQ7SmMrR6M86BVE6uJYWX
tCwPQoTf8Yz7bez5ZY4CMAKYQyLulliXG7XcJbVFsED3ugNCR/buJXb0lPBRGKlAZWwK4Fl38pcE
jJw9b99HymJjRhu6DpkykVuLQdnM2TgpH3lFEnqpQBrlibqQyfo/XZsQ/j5dOaWNtGBQLJCd4iWR
w2Y3T/8Qwoq+xitpkvqeTmCt+iirMd76CLHC9jiNjdxv1izIIivDNh9z1hh/nP8mXOYwOkzyf0UT
fNvl44ghKxAYIE1PPAF1sxCO9vMKBe2127ZnJEDm4OlWtL3IjvHK7uye8pUq3Sg9HhPYagOT0iCe
r3ea6NGDWB9k+9KXziEh+dB8sICeNRFAHq9/1Sjf3CivlUeWI3KuOIanqvRdLaSSGGbkpprUxEc6
B1pQEcbNDxnqIxleEnhAnb9yY6ZyTZwrotEySv4uY/DoLEQ9lHTPsTclNSua04HkB5G//JYUKN9t
WSwiT4UKSmqoDnqyr4bORgvgihC34Fog9LLg2JlrlSNeooNfSfq0WUa3LZxBx0KV6Qpp4ESe/Tck
0nS1OKpaK3r8qc8aXG6ER8Or7YpHODk+oxsqZFjlOKQ/Llq9WmUPM6YCGoYCCVufLS5S8iVgjlmw
j5Qab6uNZ9gdwGufgxfLCgKxza2c9o2XwAOVVkxO61Ta//4AOuFGFGOuiBrFLq5/9o46hRrMiK08
E+DVG2+vsfMqKgCq5aVXcz3tC0m3rxswn9QLfsfl8Gekm86aWNqxH595G1Xk2FFIpkdnMQBK7LhP
tZxF10pgQVln2KHoJLIGJ2uCi1Qx/v+3h4VDsp8iLwGkyb8SwZY6uT67h6KRQeKvACtPmNsRxox2
nCV6Mb5Vtj5niG1ndUfc1WxDyYdT3Fa8sCC/f17bGBbX8elc6Ji8CTnof5CpZOaxSK5pkNLVremz
59oS47EPRedfQZe7ukEKVIlsQCIcbxY8dFPFXkWtrkub2yY9nDrtyUjMCnwza8g3JR12/L4QZzHq
Rqz/j1KjZWJheSea3NWj/ae4rjnExRb/ESeL/zn7ps7Xeq4VE40MCrbZuwhJCpgGGB1J1jczQ7bW
KlbSRHpkkgWKQRUMM2GISn5FfvA9QGtKzZ+Ze8E4QZwFNC+wslSxmaJRE1L4tRnTMUBJ3Tgbxgja
AHOsfbacDR3rKDCXQ1qnFWGKQTkMjcOosh4C/0Im9+Qj1JgH1SVu0ZvlMC4r+WIRjpUbYgUlAgNP
hGkaN6oxGni/NrIZgV3T2agwf7105LM/Tnb3DQm4eipUOXPsiGu/zHgopcQ258h+oCNjA3tnt02Y
BpFUH0RoQmqCbtRr3Wlgi51JGKW5rI1sWvdLo24XrNGXHgPWXfTvoEOPevt33mcANSIOT/rEoPcD
M+IwPY0EdoLrAM7ZwCS6gy8WI8ekWCv/oM4Hp67Cgn4aMosWm/tDU/Mn4/tA0KyKPTYuug7nmD7e
WOmMRAVkYazwuNRHJFjyoWPcSdxcmOZ65WN1gSDjZKF8D8Xikir6asQnQIXvQSrJtQlOdrp7SSd/
YS7eGSxvMSgyCnTXPOelMXBnP6YGpphE19z4+4v5KeOWS6opzZwxkjHUhav9+aS/Xh4pr0RDff9u
cphgJJjHAcpO5ewJ1BZ/B13m2T9CtEAOeHWUfByHDaJAm8MBCwHMQYrgy2+4zRO2z8denyX/RL4H
jZXffg0U5FLE6FI9T2oZKWvcxvNYtA4TgXcCZe4Tq7Ivrj6MF/Y9iXaCxqJ8R9TqpnWMoYofRLua
vvbFxurRqt6u9OkYzEOa9z6KevTQgZSYi3rLa1/agedVpI0ppLuatQrRE/Y+FVXSLqaH73cYn8/D
oTKXjeMuY1W7Rdal/H/ADQuXDzmPqOdHqZ5bK6x/P49/aOqDp0tP4iFDMDcZ11HSVHMwzC2s7GQo
ypUuOIo/nulhyLSuHOs5/3kCz0MUSp2yV2vy/smdd889Azgly7JzP6IiJWvARvnFFrsbRFt2PVng
GlampSRH17zjWQbhH+ppSXKBs8lrOlrjfkACY0JFWGYATTN7KNquXuiGfqn3ea7XxNKn9UbmQAYr
LcoiwtX7yTZNpdUW7osVLrqGTn7K4WKPY00WtIngLDHi+TTQGCr9a5QNpAV0dI0YpYfNbHggPvtM
UTirCbGfTfkhLUVlq3yQ27F6Hvd+jPPA9jDSUPHOzDfZ13GJ2U6dBHt3VA35vEYPvhM/nD5sA3vD
ccdGfIRzx3n9dD4otlGyLrVuFVm40lXKR2MxwBLv6ff94veaj74zNyTF8SoXsUE/8ei2+e951ObM
K19P3ssJHJr8X1EX8QQDwYBQI3Lltl2Oq/myyoimW1BBLGGDE0UNkUlNKsHQBDlinEFWvYFLXiDc
j8FEMxU/uxj0kN1LLXtbCltNnMO+19KUXRHRoRr0mGy5aN1IKi2XJNRj6Nzr8exEbSJ0LC0/NZAZ
0LRGon4y8vACI0pdFmCx35umIGl+P2O+1Q1zZEDcdC8lgwMSGdx6KNHn6B7Jc0Bt8Fthgn5C67UC
ljubgzV+a/GS2Z1yEkXFDmWYA29pD2z4LW3oDYf567yQdzPaMUdPUGEFvCKs7Vq12T1cyq7g8Mkt
SVVWK18k5TVbVkcZEStwAD7xRL12wHqTr4Troym5G4CaPca50k7QqnzAwdng0DHrtZNgBuyOZ8dq
ZvNO1H5D+D6iP/H+ti5rjrtm5FcoIuIDZJ6KTnFqQZsF7/fR8OJ+lzetEfmLFGU0JmCq3RcQGSLH
XMsdcE+VL+ZZGks7hoJrYGCz+31dilNLYKj24vVWO6r3GJgFFJryiyhh4XzD/LL/FTmAFVZUzVo+
5GoHGC9TPXl8STzUNeovFCcZyn1/Sp3WEFV8NJAR3j8OvDZCiTLAXBxKHJYVkPsKTisM6pO0PcW5
RJeTkfctb8o669MjXPLPie3u0qkXmj2FMb5A5Frbjhs7gCjmfX3k1lLOGOkUBZRBYdUtbcQa1qZy
LFv0587DD+rf0mU5+5HS9x22CZdqh0XaB8hkjoNzisN6vGN2bE3eM+8EE6sWrQURK7np7g6Ni5uf
HdOYbGnevvbvFL/cDRtJpf17ZsghQ1IAG4/rbNeK2wd2o1AMRZWNipJKjaZpPnvbiC0SH/SL8LTF
ex/ofIFu9pfa31QnC4dNXVE12AgJ9VAD92+h0MzOqyW4ruHz5DEU9PC/j3+qKuzYNeFQdcZ1s3N2
oXgJV81Gee7AbUmWJfvX6JwSlBohIUQ8/q3r1n54YV8Q7CGc0LUMEs2W2gtrs1IFYJKr+y2j9Ouq
Dbvr62edFrPNBFOkrqjACDy08XbQ46Q4WoGfpqk/4WmnkrNx1b1T7L/4eFmks0w8Yj00ZyvLyhQ0
uaWSi0FAD96KsdHeWxMWGAEwidoIVyDOl8Kc7RoXlHxuJ6p36lNpoF977SeAIWSczJ7jDDruAgcE
yscOIOKd5WkrHNj3SyKJsOZ8puIeieAX3NmcjRdyGXSp6LUew17JckR2Hl5neIXbfrJE62/FwZOH
Qvb+aJC8EI3gUgXN8/Fj2B1+5ZKdngKTIBg49ZW8r5imVorZfsURpcDRNFdXgxbr0RKGg5gbeH6l
Xg1ZJJBJWgrMjBc6hhJY1LdzCAOPVlqkRvkiCIGdc+7uqc98HfP0887EUUwfcXqHATJAXyVN9Wct
XClp/B5Irdjqrzdb1LgSsFvgnNEK51u3d7pH9N/DGJL7xkEmky6ATdsVR0cvScws540O6y5YyVNs
mn5TOZkegUQoaa6nYqeufBWdHoVnc1SBu8K2Zvh1spNqiLWnFvkrTYpNNAf6fRx5R+c787jXmwsC
znGJhOcgVZ4G1e7h5pH4UJca6TTnUEQ7btgUsOS/3w624koXo/VhwFGlN1Nt9zf0uyq2uehPMZ1C
49uzQ9Zwbuwz17+r+sgWiArwgF5bvBCqKbIibbq2b3r3iqzYgC8F03Rle4sxasdunXOTYkwiFRDD
Kz9kIoYebGxtT0Ty+Yn5k8Oag4mPBukbwKO92FijK2/NdrmnkcmZna8YVRA5nziBRtoo1uFSTAYG
ZL0j5D/Tf4G39uzuz64S60JZ1vRlvoby7QsNJqdrgPTH2qFm19JFB25naNMla2qyJ/vErID7JDJn
FLekKcQXUK8oDyDKHS08ZMmcTgzSJqibzVzB/QE8jpXuutpmRQY2d1jT664/3v1AyIU4Wy0AuSW5
lgAb61ZSRVlyDXPPF0AQQWtnhILCZh0E3E7huBfi9j0DUMTP8uYH3l8FgF/aWjX6DORO/vlvywoI
z2FuXvEPel7V+vTFiukQPNJg/tB6QaNBSv+21SPyh1SY2KWLZnP2CzFxk1wDpOanEFj+6OqV9VKr
Hn0dDXLeR2GNLoK61/Ln5nTzVKaDiWHrTGynhQR3B+CWz7LWlFglH1bsCoWAs7BWNRNHAW+9bCDU
HtwZuUrmANR2Fe+OCD5VZqxK3GnseChIDVsoCoX9clg5OVuXMzgr6mFfUlUm/cBo90hDfpYTGsjM
z//gB0e/9N7k0gqKdWZ09dmuebPbL5E7OrrqplfCy9V7NAIQDSuVIh+wOow9KfgSRuGdYh/sl3hI
Md4lDmwN4yVGkyRUBOtjiE30wQvVWrQu6wqdLAh5rDK5s8hNsuS463b+J3FMxaNV8gnNeW8vKXNk
sVipLMy/wxfgIHwgImC0NjDtOLLVJxIOX7qpd9a4CVu+DhUt0AxX/rV1SHfnEA7cwB3I8qMIXLhW
WVxWPN714Vg3MH/ezCHz29bnEeAFLFeVImimiexLBwNEXk/bnfGhnOfO55KbYVSCn2cGiao/M5FP
NJqFj3BjFklFm64kW1VEQaXQIELAo5J55E5uxYVXqppvF6w7s94d2rqMwCkl8f5eOHlnPXTJHhTf
vcee2SF2rvb1b1TSeK9x/He36PpY9ykF9n0ZnOOy6APlbWy7eZn7YNlaqMu8Bn8KHh2zVJhm3F28
RH+V0BWao0EgPo14Jb/99GG1VABVDl4rgc8xQ9LtJ76J2agdnasqRMpOerCgQOc1bvEO6XhPdflK
wyYjUpndnRw8TZpEn/fBc/5diCtzhm+19fUF2JYX0NkVA/+GgeBgiUatql9Qjht6xQhEUCc0VVr+
wNxpGbT4kOexSI2KQv5JDx0LHr2CMc7dFKbEJT35vgCCKwmZvHJYUlg62TG3vpL2gZ9EOpsdRTwv
eBbYkWXaCtswlt3awVvu9Ksw7qdgErDzj54Iol/5tXkr7TU3cZegnkgGmxwCvipYn9uOHhmtDLMO
zmtMMcOOgszbefa/uH4zgb1DJL3TWom4rxY/hCwaFh+z5hf7kFwVd9ASEQChRoCcUl0ETNp5lryL
9Kg6PrHoUU9iwLGW9/7Mmy0LlcntrPsVIXhEXpWzUiPrJ7RKGNe1D0KyuJcE9CoqDta7nuVtrR1X
uBGbqLE5vU9odn+gZNdU6rIuewxUQWiuzD/q9fpEzIp5IvgOdTLkhNcdIn6qN1gJkfoVLL+bM2jY
YxlF48tY4VRRphp3l3XSrGSIjwFNOS3XZAf1DxIZxZrdmCnsoZqnH8YROxlQ4hIhTagMur27y/ui
rnM6YQejFPNNAA/LaokKy8jmW0dPxoovkXwTq7zyhdOXjnk9m9YynpmPzt4HmxYBddNgL8Pcz17+
Tpp4Gja0N3AODB0J3DYF7ZQN8hhJGbk4bLJgwSr1keCcE3BLIrMQymHfRS9wy9pu9zlXl/tUZuU9
3vl4BWe64/NJ2uwqGIR9ZXShkGyqsu3xwwcJzOBxms4Qj/77DG4x/gz7Fa3eeDBU3Du8Gc8rfvnR
CZyBIWWXmBxhcmVK4YhJUGLJ9kVRozqa6dteJaqYvh5TtZno7EGMvH8lW4iZmWruJDU0WQsWyUKQ
R760sMey3de58jSPWUyzm2ug/yzSvebrTw/rGHVo1n+xuegXjBHr2i0CNAQH87SDF3JPTeSGokrs
vzwAAkyROYjilf/mJgxuMu+i36O21srDhOoBcAMezCk00M//e0y4OT70sZaXxB7iktgXwcejOB6H
RA9+3sKeskIpmiFnQP1Pk8Iz8JmLxmK+cIrsS8QfmIj/rQQCHm6Dj5JOs0POvN47I4OU4iyK7DD1
UALbI6OGrXbxCPJV2hjHkOIP5iVbZntmNRmwxYur59IcbAQ105gCzVQjBlmky7quQVrls+x09qjK
KHbhf/sAaboX29bJAkQ3FqnKPKDBiUGMAlOed78dju1kzjS8O9Pv+jW2uP1+hySODjsGyqw1yfhD
lRFoYhptoQvIYU7es/Fo3VUgGUgBFtubMdyhf6/siQmbWBmO/HXvcUYynmc46n2bjM+hs4ie3W0Z
RUMqRari6ChUi5nVg4DDE9W5BbJ2isebn6APmYqqnpY6B7cBC3QJ1A7vWJ7enn2FoMYadObRJ0Pg
Ht/EW1bDeFzt815atW1W8H0i5MFBLb9YYC8VOLR7HKFEFJeckZyOHtpZY1kbaSEhNhLlX5LwkJWj
s7Q13UF5DkQMM0C+fFWbnmgdWG2NShdidhGdDv7YzNkfCCX4tp0zah+QHi94t5BhfkIvK2EfmURI
voTHzSRjKnxfLvLE3mwkgNfurxCZ++Q/X8MhAMleq6FIwHaOQGnjmZ5h30ntHGnV0k5StUZ4Fpbf
vR2mh0uv4PLwD1pBLiRsC3FxSh1n01q8MyTUKGivMPziolB8hU3BN26vSgicvwnGx4C9ZSKCv7q9
zoFonK/q3rkUU0LetVf1xa9RrY7rQ5dsomks7IMmr4h1yf2o3L4vzXak/vPk867OBB4ZVNTYYtDn
qeW0O2bFTQiIRddkIfuHfYeDuIG4LqaMl97LjkNkfaBW5Sxb0Sh1+aARb8wrg5IyWD+trZMhAkJq
mSSCMdw/JLmj1tooSYp83MJ2yexacR3a4drhChf+/Dzg17OAZL4SWbat4zOApIIqPVVqhZjrrXtF
KrUGFV68mxa9dG5PQqhQ/WE2qq1aqZCOIhbpxByhzDCpeSQwpRhSRgixixWlJhqSHek+c8/NPKgW
n90d0JonyXMCvVUgtSwHHyG1pU+apio7df4HYVGQWAVcSohYn/fiD4VssFouhsXz9VCAA7AiqahW
C2HfGgaCMxhnjmTZEX2XABeFFb4yGoPXAysXG0jF2iNRGA+7uWm043I/aFUZPpKEq92Sad9xj8qv
K6Itvz46HFsR6oWAgW2IR+EcHGXSbmzXpZ9ddQla38uwtwSPYm9pPk4p+NCpzo/ei3C6+hs2bapq
iM9yx9kC1A4mrf2R4xH2WRF6Yymef7T2YVG2FoKVpgRc1HMteq1hfmqTiFuRzcPLAzCptC7zDv4Y
uj4QXovmNB6JArhPXsHfnZhgDV99W7Rqu9nrBixzIdO7LLvSbNmTCHqBhdFdsUOazeH+xyx/5x7T
/ui7bBE/RD4iIHGfOAE+tXpSQsHNvcG3sjCfmkyeSth//bwyZGeojPn6sCFl06EVTEnLcZD9xYUk
Cnr57TRZv+TYvgVjbB+BgveIJ0G7hHp/sQaEQVB4tXm1cZgw6XpWFWvqjneHFbauPQwd2rvweKaq
2x+ndUPOKR7b3Y0xjV3/10HPlscKOM0UiAr2KjcBVsMumsy76pfacOzBjnOeY8XuurWH0+ilXE33
pQFKz9np3jMHG+JAg+8K8EIVQ+YCUoN7/y48OwsvI6fHTVttoHxHsz1AlEpDZIJGCyAyrQv1KdEH
bmKarjyUoEBcqAmeyNpjyzYMRg4Ao/0JPghUI8Ufvw+ARkGOnZDQxs0gKYXYbjRteU7cDQeJmYUd
hFliLSynU5zV4sUfrSpqImYDUTDNNXdyrgF6hKj9kRFu4Y2abwfsfGX5ELunDCEKAdO3qO8r9m8y
qU6/HRlTFJlz5kr4SlvOul56VRPauYyJd/vYj95hsbcneG5Hj9PAKDVZPwFZqcLeqe7A9GOLD1f2
YOfDclqaHGC9VU+Rx6kkCeC7vf/WVjWSVwUxOhNv0kek41veow+2wj8rnj09YPH0egMhoYKBVDTc
LqPClVvXrsc8MzR+NFG9L7TA8FobGAj9riX3ca4ud42xQ/n62CHAntVFLyPM3DoPIlugXTR7ulAK
YvjyG+48Cx9jOVY403oOZ588+Q7RzSlxbGp1PCwaylMTK7egvHs4P1haUQCrNdBWAE3PU5Dw/d3S
QCjBUkqrWFVKXccNO6OPyMYA26nOXb9PSLWk1YIozzCb6Z1g/CJUAYCcD0lkskckLRImVjYBF+Tn
KcVzNWFKoSNP53EzvfwZ/pG8aI1UNuBgYHKpLNuX+GUVC6YDL8hgEgQBGOz7kARmLPKvz605vXgE
ofFbaE/obPBKCKyjPacGCwW0038iwo9W3W8iNb1axd0/hj2WKT/rz0v3ISENdezWJu147H7lUXH7
54YxfIJ9t5yGKrT+XFLwKUaoihOjhuhePNfsFK2V+ee1VWDJchljdBUvNtmLVQkQzN8YEW/qiE30
flNxRPO7WzGqjTT+AfDVtLaCy1g3kmn69gu9HfC2C+qQDQPFgqu6uwFrihsTAuR4KWowVHC5D33n
ZQ8gO3d7uxpD08br7asMUAg5ZGVLNLPhSTnkBumfJaA/i2k4F70u1gAr0x/VNqvcCIWX11YGEF9f
lIGMhdPpyfdu20DtCCHFV+Teu8AxTi9VnHsAg/CHJFbsf1evkGQM0drNuWItInBbQvRWlmGo1y7b
0Zo/qrKdRVjcrX7svd613LimeTw3aJo4Vpnj0L16UBue0odAttzPFyPkXzNGBk+AZDaGag/Cy7i5
KXJG6sYe1sthmruwPeO0wpp1ZNKSv0UwZ4x/ZasW3Q4dsJUvFljv1rTD8+KEucRj4DsSvjdw/IZI
jcgt8qqr4T/gSeTvvXgLPRsm3b1q8ETrCpbB99uabiv5nVDQMN3+mh1yE7l+Z9KwLYEBYWf3OP9C
FY4MK9pI/3cs5fZq8BkfFct1LdO8w1s6DOhhPPUxxYCHKZljq6e4huokkCiHDwIUstCI7gvPHzVS
3cQfWDCYGF/S4Nt01HQ3Y6U/pooVf2p0AkHZ+U+vTLDlH1gJaWQ8l1DQ+H2Ja5rIjtf/DiRtKrPl
y4rhAX7/Q3lVJo3m1M+ShFMbJSY4ut/7BHQx08ILZRXCw75imMWz3VKJSNsGEhck3hDOEGOs9XWm
D0BuxmbJP0QTHtbFI9lzVzxhB/G1eG3TtrayEH/9GwziRiNSnmL77vhIHKEXStsG9sg9y9NponFh
iEVX5Z8XCHzHxgZb5Zx8qbLFw1LEiS9/nU2A8DGLA+f+vtBCGEERx0otUM1j1FjFogKwkAj6TcYH
PUr5bYItlRkwQD3U3bC3NRSATEnTfe8L3wYN8VomACJM9TCwm3HqpPeptNW9MEU+XBDCcKgHdaLk
Y4+M0brBE6OMASZbA2aAVp6vi6+DFH34l7q5FPz5Y762iqiySU3edadE7N96HhpI2VBiZyBW7zV0
MPxyYRi3u/ED8s+599pm3zDZcSTl4l70q84KWz/KOVm9o/fDP1gpr1QLo1XRli3D1HdAwLisM+KX
henn+trQKhuLVUd9uDRYVuS5WnOMfFqJLu6QIAh2t63aiL2oYDHKR4ubpnk57TgGUjqCGobkiAsd
PCi+0Uwx4HScp9I79jd5o9qZEVA+wimz/8Gsm78iVgvG0WpzYsndluXyOamrqKhShyYWJ7CxC+lI
bjNdKBfYoD7SDJrA9P7gkcwQSPmcHb3qfKeDoJJ+v22BKFwJR/pER6skLIHXWsyATMv1eutSmh5s
HCGsECkeE2ArgrF0lHR834rovWZ6uu1aq7ip2VjhhSdF0DJgJXCIFoGvhNQjVOmDZSQksl+/V0i5
2+Y04weVusss9PrmBHDXXunz8YDbBWxRLBetozJ/8d1BUWl05EdEDWdQex75LABkDWjQbnamsvoD
7FIwQZMaIJwkbE25Gas7BKMwAK4+AfFSLuO9PZENfpfHEyY4BZsRm4j7pDiJbrweBTgjYX8OHfJ2
q+mkfMyX2DL2Dt0ulrv7o0VfSiAG8EP71m1UFmwQVeSJqjYwj0CMGfJNWq+i2DRdlYDN9krDvfKD
9krvSqgBSy5U0W3dksYGC2LOK1/K6iR2CIQeflyrK1ZY0qYZQ7o9076Je4Kx0BfGqyZaH6QIwGEP
rGkyrSZIWl2ZoPhSqFc6OEdSSpILrrWR9Y//+OPNssDZFzPgDeRc7RIkkeXiEUjvHrTVSncPWNmd
32so87y7+YfCjtIeHiXQdVZeymG0lfGzlR1GTcA+KqWpjIfCy2VtsKatcaQderDRIcTlK5RkpgBj
ljAtB1x9EPgDE/MyP3+RPYP+ZubT5qi4/6S4AU1S7RgIe3iDjC979clo2wto5FfssjUMDjd04LuB
YzGq52T75PkSd3Mo4nFrbl6Qqc3/R6QZg9885ZPFAH2PGswL5gRm2uz4n3ERdpYakuwW9CpHUMHJ
K730d1R4bq7S2cnhv78MHi8k1I18FIAG74tsONTJ5cw/370pANOLByg17GvpHFCrysTlZc5PSJkC
66zBKga0esC+DGClSA8gwkNVVbgJP5Q4mErIaBKB+4j1gV+eeaUBIhTCakZwHnbh4+FTCjGEEzQH
kYVjbdQlbuAIAry/hXZ4QESEGII4TDG/uOWHFwTmTFEXwmYP65uiSawbFDNNRWP18EoarEA3MdEG
mI6zRtmOyYYH9ui9sGV85FYiM1ETdLhtVzV0qNhW39ors/SPAVyGrMnJoz8Zy0699BiVpFgJJDBr
P8k/qRvoivvY5RZqMXUyufksk3knHX0XlAa2DO6CLOmlC+RLGZIDptkdM+E+IvspuI5Rjn5aCr16
m0DmKQHUOcEWuUF9uQWAazcsMZPOvm0Ztg/NtyuR7cCfYQhRFE+XaxxduBu4GugO2BBzPnU8T/7Z
lvurJ2pAh7A89t2TBy9DXLpt7GHeHO3hCWFfbKLEDsCgX0bXpjbwqQ+pMIoa5ndgY4BASO570maw
5d3Q+U2LGcCNFETZIedf5MEm/y7UvzTHAouhUuBxLcihTIs5qhQHAkNF++6BwZiQ3ADLqY9bRX/I
lGj+w6ouVsXGfmyTeloD2U+Dk0yLJB3ec9veDNNx9QeqMAvDXfWsYxbHXF64zglr8qHAtUsegN//
ADeBbUGKO7vfRVGQZMvG54MZ/QHwaGJY5uYw9G9DLFaVD/pICF9nQj7pQ1MBqPfj7dEbGUCCUsIT
ezqacRMdROgPEi/3FUF/BKNokUWHw7oCYcPlnXmGwdpz5viTtXt554D1Zn+krlH3ffa9X1oJJiYe
33p/XMGWHohNb8pTFYqXxe15+p/S58Av7oBjoJE24wEeRp9QPYhwCNUU8FrM7ilD/Q97LvGMdNBQ
wfQ033zbcgG6wcKjvfHNreOTquUvCy1E41HHMwIZpfE/PFUBMO4jVBmjZbj/jDf1+DjVMRB6c2+Q
ebN5qALo0r1AGJF1GAtkpDjF0fpSZj2CNcvDUrZRfk1KY/4nGcj1fliz5aihfnS37WHkb1oJKA/x
o+aCQgjlahxItHbNbU5tmd4/Jw1ybzktw0zXCUS5yF5FkP7L75eA8JPtwOTGY55biTGGXKW2IX8N
+I8rjWvpS0yx1XNo7pbt8z3Ottm0Q1b0eHH5jBsUtAYW65CS/4KUL815nCs2jHMRvFinh0kmhIDR
h8M5VLvxVlabHOabxa1LNw4eHB+BmnOeEhUbVy7EIeKyq56XF3+UWQllltLnKa2CqZVM02NXb0NJ
/cOaYFT9yX04zdNSxLa0qnLOyLKyxN/PDO6E0OYZJzkmjQsF3rfyyiK+WXO597yMz8NtFyqqIe1w
HFI7+dRDlp7DqloxofPXbPZa7SNPwP0JhSdSywLmckRwsudUJnkwwBMqeAidaXLKtI80i/qUQi06
R+38pdWL2CfoC0c95EkcAqqlDDOYRGx+G9h/xnFPpaRDxZ4EqYg0nFb9dOwm3AmHkGj//swj1hSL
HAmkii8vl/CnH4ENE+lBG7Fs2K9ANApO1rex0krRZlBuu/ndb6uS8QP0DpykiIiZlrdsEkc9R6Ws
gCYedljeZaZdr2dudsGYZ3I77gUrEAUF3r4eNUPwe0oJCbY6nVAdEbBoBFhYVDcrGMhysH3QysgN
udhSOwCAccNoXQYMoPeTNF1p5QoMFjYsU3V2hU2iybH7k70nxaCr2SUu8S0Plu0nrG1BMHHMiCx+
QeR5JenTH3yJuPPyRmo9/A/ITr0zlxwaYoDuUJ7jaCHLNzLxPq/big3JvCzdx5xIQ7jOgZmo2ioD
RmGiQIT3ex33MhNjzgc0NWFU308/0sZiVMg/4DtIl11CMIZwW5rveM9cZLDe3kgsuK4sHr77oB3a
JpfPBEy+PRsNZ/E/zSKt6XdD+k9jJxxoQyMaH7NQz+L/Q9nN3YMaXtj3whUbNY6Ma8hHfGD7bNaY
v3nuV4iY4+1fU893AZO1GHqKoOl0m4thVc/anzbNvEgzReIfMRi+1gFWF1tPwZMqXgmVxDvqPz1R
FtbKcigQ+SU+kVz1u88Bwgs6FbFdO2VxFwX2jfKDytl6XJmOCU8jrfc8aBUKqXVbmnx2twq//5tu
6eGzwNGF8j9e//9zuZeoji+zKCffxl2ulq8zP2UqJVijJYzarF/c/3SHL+LnCrltTc+k/B663GQP
2Rr+PlsaOAnIiQDPwBqjTIJ2qfwscLeprPonbmA0rVRjwy9EGuhKHGG74TRgM3iiBgRrM4aU+Dms
0ncV+F1Ac0ljnbhgzUQH5ukcGyr8u+VMAPSWUHiWB17f1KaJO3vOrPM4iT/7OhSWhjadxOFt8AE7
tvABqOKoHbU41xS/Q1yRIC8YkxDDYp2Xtq1IBMHhTKeQHo8cTlvi+Dgc1xYYIs/gG2ooNrLb9Ijt
WTDLMfHrIxE3ZOpCPqWWzXvd+mwsfMh9HBmaz4RhueQeRWyIOwOdSaJllNRXeu/QXUMyMfBiCu9S
lwxdY/230dC+UP7aZ/gxv8AzdE8lcJFcsypeKxlcQBUD901CeMGFFwjYlmLejAlpoRCbknI75imV
e1ZGhIPIWJNC0meyfAbsYEs48jES1zHzS9RZ0XeqyTqU4O8oJtRJ99/gTqISm5jzM5NN6ItVUajU
SIyULeSBYnUq6GsJP6AgyweO9RGYX100qASHSx09jobqnE4f61OewmZDHO3n9g4qrDJHc/H3mQPQ
GMFWi7r6eWnpwrKihtePxRB9eoCl7E6DlJZj/Sun5+iKWrrZ28CGiVs4QBcuENOHhf/2WC2RXe8V
ypRGNCahgqUf8pDFngbKXmUAoK/XIkIdcbOLxKZ+BSPAQYGfKvpiDsWr1baA3eaJLwCnAw5/Sd44
EfOXyoYTQwddL/rmQHgbyA5e+CeTaRRWUCnk7z8qYBv2bTTuDitF9w7a4+Iw8fV+yKzX2ZQcWuTA
G9s7pqQO1F/S+u6UwMFe47x69FtJAPg8pH0yk4BEvJIRYsJtjlByKTxXQo5OGIHYtA+tLAbjSnwI
DqNQc3NOFDKVzX4VZ7Qt4CcmHP2hutRJTjPQ2ZUAw8GU6tQRTRkUKthUn0XOBWI7wG3QCb7Hcb3f
L+FlzNYMerVprkJnf1D8KT9ee2HAEsydBawaHzyiLDt8bilGJmlaLZjwKH0VhAEUdNs/8JjkA9AO
dgAjhvYDT0NuiicbUjt7YgaldH+ycJ2+W5r2be0U2949pU9yOAFvSV4Fj44/qa0zAxPoaABs8QsL
kdTp0m1824hUrcprmdWS1fOXV43JnuuNUtHtKasbb8TwZPvYlUBUgsp9fXWm0kwp5Pbs1BmirhJj
zrIqMxIE1ucwd/yKMWUDsx1dxNFfRbE3at2Y5v3WJKFkPPjtxcLgGvxreZ+Xv0a4vdFUihMhIK12
2mRD+AiQyNZU+AQpdweSI2DYm3/5omo6KwM9KNXL/Vu1c3NSx2Cuj6BLNcNU+KnxNEB750aKf0qf
9yyDFp5suhwm/McdBv/3di/ZBrY/+CCyjjiT6GRnW7G/TaCtfdLKeuCfYNeEczqsXM+6FHNAIBw6
7plIy2zMQ0Mwv0DxFll8MYo+tu1KQU5G99a9GlYC2yYZbxH5Db2gMw1oGUDQsXU+UJcjsFpVXQIq
kiDpb69T1KoZXGXz5F4JRvz0TqUMBOiGr3Z/1CuXoXO1Vs4w603yF+k7wZHpt/IrRU3f1fBaHhpr
XgWWWOUKzf4wAXfqCISdnxOPgZjzzK0zSPPMQWJEb+0Tm6D3/F99EsLs3tbRwIJsnC2WHHqaQAvO
GQzGuO+4q1klgPkqIArZBih1qg0EC/AhMAynkHEYz3PmJ9P7Uhd4uqEz2i34q40rTkw/iB6svl0b
70A/WQidnhMFCqwFHP9KuGqc6EDSZToVJGXP6R8lAq3Rj/3OD9XVVEkO5HOBbwtDuPHN0af4duVw
t9o6Npl2iZqhzilldD//Wboa5KSlmUCVoA2KFK15F0JUDHNZcVUENHok2fwI762/lklOnzn68wxJ
RvLTX5t8ZCnhpeUSqcEcCo3rGabkCAgZb7+veCm6Km+cX/bXWqtp+FPFlYZw31A55uhiEyDNXAGM
D0YzQcLY4NdwzsXqLdVEpPn7sODi5JZWkMDRhAn2XamjBJ7gYwV3y6JWsykb0SbPvApMBPm1bis9
7dq3XYsDNy1Z0Zckt++nLeSPSkWuJ9HNYY539P6WtHFjzNguf3S4MCb/a8bVTCsOGhqMXQguMqcw
W/6itD5x6Z91FE+Qaakyy9s9ea6jiS47ABFaU/L2+2bsykBceXmHfD9rY1DzL+CYPT5LXUwvRWMN
qfgsIfyf5i1u+1QEQ19pfoGrgvGHsp58ZuADukgHnPskIuTgLziOhMdptvdMnfAWFlm8kUNx13rP
epxUkItgd2sRQSyEHgwFaJGrXJNNfWHA/gwMgI/eSxJwTxrFCvFPjodUNogQ5BpnxwD/sQFXmSYk
DkAarUAjjivlgxut7i1d+VOk8/qNBPj+LZhdkQrNRssf7sOvZe+x6QvXFacmMPyILWtq0LTbuNC5
Um/7HrngWpusxGACNvdtAJ7b8dE8n6FnUVgnmBFGyIWyq0bkc7A8xGetuEra4CDlqMeqZJ6fHcHc
cQslbNxnioY/+/cxR7xJHGE8wEEjtPa344tllg3avTlP9s/lDOlvFDx4JMXHwq3wSzgC+OIZOR+J
v8PfjCqOojBp9n/OYJZ8GUf0NNvKwyJ4Ce/d6QMirmJTFJl4EAwZnbXg3EhBCa4Oac/XVsrN+AUV
fRd9og6GFMH3jQoSnahCky3q1IPVJhaic8xAfvx3ibiYPMjDjMRe/b0TLSScSmAm9+ZaxadR1FtU
jNpckwL9zkdA5BsKNIQGokf1huaH5WVk1zPOh/yupDdLGMiGSFv3eUn7LTJYc6wQAUhdwUWMA+AH
+FnXhSOvvlsbQ8mbCry1b9o3oCavaDnLmxpStK2Hcs9o/nmg6cl+Q67YgZxMGAL9+moxvZL3O1rc
qhLr/Y3+AwYs1npF3SFrehqfmx2CSIFDIvIv2uzaNh4PkqqSlBFsVNEIzsQemd117zS5OHlpTJ0k
9QnQFYGycodbPyGHwLMA2S01EY6CDP64tXiXfSS3F/Lv0eKCJCdhSEXQBQzNzerVYjAxdn+LbxFX
/mKI9ALNP9HFcH12Pmm3tpdUWG2CCda3dyYOTwDkftfTeD/Kg3lZN6iJawo68E0VZZqLM7EOVMqv
YmtC1Fw+soMWtsSzIrBWIonEOLrB9FO6F8XUF1McJcOm6J1fzLcAob5y0TgZfJLbM0qBHRaMdSNK
2nB/7rdVZanwvyOEukeaSIHanJNyuNe9tO3Onq69l0uw8TvbOHYSRK0NEiYQnwGm9/sRF4UP0i37
ooJOflaL0QQrJOZB3OSCZ5o3iIZpKHGtA9JofEkEt0zp2+ICPCz72dmJYIci9fd0Cb58IrkPAVUX
WXijGbOdUHzLD1+qwZoIIns0Y7vsh4lG1Bd4Lb/YwWNFtrbEZHJRV4KZfn8Vap+0sQLfMhIm4FRp
m231JUwMlUejTFiOuSuwzBVbW1a4N83601zC+OPLglYIVmoRcEhfoH+62ioBnjCGMi9tbXUbJDFb
JMBTxUYBkap3Ox8v+BgnTnxboaLbf1c1xmn7gYnWu1OyXy59d61f7hrUfB34A926xtQu8UvVXc+h
aUMknlbIQ0NIVtnyct/iknYTy7s3RWJaZ5ubrem6vrs5GEBq2n5+9C1DwaNcPTKeVgrPsYdCNrtO
5Sovr9B/xltPIWNzQFyCTUKq+j00TkiMLzO7WvDeCtAWp/Tlcw95QfGRYOf5jDasmlgdGy8jVk5u
UxkODdBTh46sihd1RPe57NixdRwVtqXrn7ixGbcUSbNwL5KphMw6hJXvKT8hvHPf5WmFJvPHO02d
es+O9HpBA4ZZ2GzG8aPAetHZBppysYmTXQW6RMQrchAEoUhJ3Z6stIKLa205MIJ6bDLZwYb3U0KO
Miw47ZN0Ead7Sw4/+lTg8TSH8i9geVCo4qazuo25GU4oRJbAa90E7WOjQUVV3z4e2Lt+wYby6MBy
frTxvK410AXpW9/Mmlzg6XLQSOwU5WLDQ16SLn7X+XdIlNuRwnbZsieTYTHvBAWtCHGDH/3BqCXM
RyPcntYeiNeS9AdGEAU7KIrkATkc+XRY/aV99L0hv+6xrTF20/GFyv1ycXyqbqp4o9JsCqUgJdJn
MFapseNTjfBg9QOQIK9xUQho6QAc07DjoV3rqc6pPKdzNule3pw3RczJrTGpRf5L9gCeQSjCBTMG
eUuVMPUomvD+eYKiEsBtH9ftkpPgTI0jw6Oqg21KH1cOu3YspCbpFmr5tuacmwtOC0wJW0odM6cG
sk0HfGisTHNbiImb9jf8vyJ5dMct8ySR7hY6Xr0NibpP1QeAIdk36jEl101Kab0VuTXtVXj6bxsy
m727es2Jk6c6mrqxAoih7mpmk61jg/sSzcXrQi2asLIL6PZ2GLCCxpY7PR6UdZyutVBKFW+xhiBb
Osj4XfdMxwS0R/+Uw71urtOzzrV0Dh76cCvZfhuPy00i2B0oBvqZgjf5TOdxJSrY/WIs6/g8Gp4x
UOSUBOOzhXJ6JW7NrryG+iURMpAxYJVyOOB1D1C59TlZHxslegu24/KuXTz3Y+/dV7HeK1qO4+zh
MEOabIR/5p4BBaFWSyL+WZ11gA+Wtnxt8BnXaQ7ydrfBLf4EEU1f8zLY8pTLBwbTT8Vvr/WvEpm6
vEeImKvQnz/lYqyOHmhwcgnCaYIGE5yLOs4xemf4RT3NXBhi0+kWOEcQSr82Sgf1DQuVesqFK+oI
xcUi88TMgvHOSxD9NK01YDMft3djQZlX8F6Nj/J10OVgjujLE2Bubpe2G7ca/Ke3rUV+OqnWyc2w
IQk+8IF+YYyFh+mBghg79AFoo5K9hOYOFAP2zi7t3S+I9LR43aAVOPTTo4hIppFQDjtQWkI2teyb
G4+qtRj8njWqtX6H2zfjQnIrm7+blLWdsoEgFl2QFrpKIi2O5Pmu8V+1Ly5TIj1Pb+0HgLuVcP8x
JSNpauzF3hj30USQnoHQZXcQEjpuhmelGS/xpdMx2+4KzBUrN39AbZpxVBUrVsp/qDwma3SgLgko
v7I5WlqDlKS8z92K+/PCpzVc1d88oFcgIo8lYUaUU9Dn8t6W+MD7ksTtnu/6U41GrimNmewpViEc
/pBfpgQbSSavFfR8MzlrsbOJY04CHDeTCHyoB28C7UkCiFfTQ+XZyhT9owfyWPp0tvWVs/XnjafK
CgrhQUlQUoLPE2hbAEPkTBVPKI0G3L+lSKAMONomHwm2vPSztFyawfv+fYI9xwlW58t8//csLmg1
KkJMjGZzs/8RSDNxymndV1Y61ZDLFNpHVcvX420jGI3tthu0dYZgTgh0WfYI0Wzn0f9HlTqsQ0Mr
8Zzd1bgpRA99SiTMqYjIjheheXb4vse0l575/rLtv0BMWe0GsPXAZ7K6O1tGPX6LSjlGOnJIUiVN
OFwurc/z5B9Ll+vUhihwiE0W2oH7wj37aRzH+FU2+r+lo96IYxA+8JA2yukrr6M8LXVTTo4jGJUW
3/L2wREexKEbqjM5pPNega83Zy1YPbwd3dEGSvnSCn9VIk/hgL8SsS7Y5Y92IlcGkx4KJkOuSwgr
lVxLZE+aGc7qSekT4KqFx5JIQC+qx0m/glULX3+60wEdi7WHa9QZmX7NLv4OcS/DxCkCI3xx+bu5
YCm3TIwmyFEOaWOBNulZuB7aCw7TWaes0cJBgr5L9PkJRepVFG/kywtbHs3JAFXWoczvQ159mI8J
O2aLQV0IhS6lidNM/ceIPwRp+gtOZWfdSBMedIetIsjOG0KGK+sSgodmbsQ+vqcLWlH9l7kecR9m
+GZv6+Z3DDZcq1KU+hLTiB3tbzfv354/pS10IBSivD1UmEDSk5vO7lEhcUIp+3xO4e0HL8KJBM59
NJh5NmjZ9lRfvEi/s85stc4itwK7InqmShIB4DStY3C+Ev2Hg/7nXgAXwOrICuEVRwE7AxQL1XXG
JIlUTrKtHy0g3feeQVYU8g+D1bdC5J/eban2+3zx1Rx3ZrX0V65vRbOaWZGLEbP0T2miOUqaR1Fz
RARCeb2eDZRuqIJBD0NtJ/Z1ujdpoS+ifeqwGgKpTKWeXFOm2ENZ6ljS1/z+aElRvMwMAS8XjFfC
6vPX/kp1TIN/6l6zFSnYze8uh8QE7SPYLooc/U1zNM3sE1Toy8vrLz9GgPXYhkNbpIq2ye69HznL
eX4A7HYWlL0L2onxDyYj5ZlvNSQT9rYCQRd8c4yDY+cy9EipFrg2ma2KA4qK8jTdwdrtO6nwrrXQ
kedrHv9/AlNVL0XW6travU28AkPARm64xyPG726gcdAPDu88CCMaNLm/lO8baHZmJWTYgzUUGPnw
6TBMW/1o9Rfb054fxCnH+6eWoRXGe8xijcJ3ddYppc1MnUUJa7/5h9i+s+bFl5fL/VnADKm7by41
2CHCq6DYIFNWahC0jTBiTlurlPI9DFQ02HB13k4ltCDHdzykpJUtc7xeROy1FT2qxVEDEJO2ssxq
KvOnbD+UGBibTgOJMF7Bkxp+U8faNez25KFTy0lMAUjTlFLreDXV9YxpVr9JnbeK/UDUNLLLBT2/
w31hUIXT+2iaLchOePaAnHqCLtvmvxS2mYA+000HOQWfQ6FhxywynI6FyZA4ohfQOa6n7sylYQYI
f1Yd+UmRAqJfDn0Co8YvVtfrNeoQeh961iz9zTfRo78gkRHEO4H7ti+m5mBxN4Cu9YRbbkPjpczW
46UREelge7v9Gqgv8tC9cblx6zQc4XP9NaPCCpd5KsI1tCnsYWRux1PgybOB65NCVefUI1m3KKfQ
nrF80d+OD2ZmnHifigxhDVANdSKBJ4F4XZwQxH4APW3NgcgwlfRWz5XzkId/2QxyV8x7NAV5TVAd
mdK9COf5MYJjP8Vit7bLaRTbhSvaNHkZMgkMp5Xw2uwtFnPfqleHUKG9mzoEGKzg8N/9RjwPfn0s
V+eBlBKW5T/CNzf5TFZU5cHEXNKnoN4LutanwWKELCGWLZXTIfppiba5fbDd+jDaIg8OU3Wli5yW
M++A12TEKu2AuuawVbgnshdWNMVLvaMrSKJR10/rOTOTuOJzQy3LCkWtGN3ptSxTK//aNuWTiJlW
47xEmBGLCv9wU33ogQF8wn3JdJcrOHihO8toQsjeg/2qMFXa95jPBY/XYxudsmYFEdYAkKmoyLuZ
ryi37GGQk8yz1xSIxUynVC+V4yIOnyq5eK5Wz1WSshjqMWG3VsBce0taG70wS3kZIq30e+6y2x/e
7vAW/IBWmvCjDKzNm1qd7CWULPkoztFUTlHm/42P+UisrpK78sZ3PqJ/ax6Te4sFoHQG4Y/q5Ihd
MJChMbTsAJDoHdOss36KbHQzHImUWmedeN4EE/nwgYZZMQXBhYF19SJWQupb7bB+sfKXO1Hr4RNW
BFu6BXumvwvh+DyTi0TI/ETXvCZsKIUjWiiw+r+p79yygRhvsOQCDFhiXVM4+jIudoyQfKV1uJFL
Cu++T6qzBn2ra4cgHJpyVQorNA7QRVigepdpjDVwwHR9YFY7grF4/mA9rgPbngW6GF2oNBRurkbA
+UlnU0eWfa6cEvKfiy/I30XlokX/+zlRlihdCqFBYNrple0gY0FmWoqMR18gjCItuDfhTkaBlRWM
vm4SG4vt/pIXJpbrEVyR06hcb8NTgarrN6NBAuCYzX1ZXe4FngzPLnS56PvppYdBQ7sHn6tjFbBi
8FJTE41FYJd3Oy8KHVYZPOuYgph+UgBuE2a562j+r5HChXr/Nn1ShECvnNdnRig+4G53b6qzOns2
Oebce2T38tJogJRB1T6spdBUwelSEsf7CGvFjFaVkr8edoenM2FYnVREk1iJUxlKvN+XOPSD3Bo4
pHTxCRGBEa1rvCfM0vf9bMZdSPiMi3+77xKFUSa7eZI2nciS+VgXxrwfh0qpVwvAEjb3N3TGytiU
kj1H4uN3CfzaMxaSoZNU/9/52AI7rLPy6IaU1WOzalG7zuiBb4j8BbhYfvwBNqD8J2qGfQLDQgM+
PrAX6P559yaVceLRYNdS3UX0BttqRSZPxVmtAHsdiE5VwpKAJ/CBhjD2Spbb6DKYqjm06Pv4gf3f
5UU8tpn3C/KrnjcHtsBeVoB1aemg2lZfuHU7t4M3W+tYHPE3a9uUqYQ9Ngio+GT/c05AzoA6RRsp
SdMkBBnihrWFb9iQ5kY8z4eCSC06zW7pmNp0EX0e47c2h8ve+Q1yzrGJDOPkPac1Qy2x6WyHHsxP
fO5J6G74hk7iR11tEfa+qyiDFzGMPxGPBN3mIBJ7vPwsO7e3F2Vob/WpI4CvUSYbVE2k3trgfK2N
q4VrO8H8/Ze8kwuWc/pF084+cEFI3ZsMB7i/uqEMASX7xqDNcKQSvhJdlcfMtb8+j6WCYefbmmGh
218FKOUe9NsOAczU/uMwIMKQPEqedcxlknWWNtiXVy+TzvCpH/i7nGuXyx5oqTCIe/NPBF5FQk5/
t/GpgU6v/bqqY+WCoIinWT+W4OjwFKVcSdfMPAEnQOfeRmpNyO4kbL8VpHnsYnvbtpRF60L9KWQT
rzM2UZkfh+/e4wKoiP9KWPKILs2hfAh2c8BQ4zvUyO6OS6GwTPIznsN+SMIc6SPLMmC4SMBkEHIE
4EMKburMHueN0YsjrJ87+vDmIQg5XrCEbDAr207NGCSLdioVyBJvXtc9UBOhBvfI7uX2RFvNo0fZ
Si/h7kSHau9UBI5KrLKWlXR3TGZdB1vH+aNDZqrAuCUnzMH4u5xNvjbQsJr8CaV7PoU67P5ezycT
uzTmKgea8MsglybiLSaSOJ8JCawQ5Ujwmzsc7Vq5t+yG2h5V+2xurpp8pBjrEggbIYg1U2li5KIP
gxf5okr80Ty4KsxVje9kbC3ZNmkcuzatLGtb8RVP4D5wMms4tdcEIKm33nBG0yDr8V/7PgK9wJ3v
3RB3FCpq8bfQCoL9W+T+naFUM75Gp4OKZgrT7T+VqqXIyoWr9X+KUTVvdycOuHskeHDgLyr+rbgL
8QUoLJovH9q3i6LRb8kuQElHKc020eEynMH1AqtvOiF5GxgoRnBhvAljExKBRkRN98IcmCpljzSX
b7tdme/HYVNdB4rlbLBMNbS91W1HHtFrFGQviqJYiKXATWuxG8wvCS4ABLcTQjGwc7LvsQIhsdAi
fqGTMXPkcYnse1ZQXM1zuWIU7MFGoxn63hEt++wYhs3nntiXUS/6uxgItle5oAhzxo0LPckEra/D
eCh94KJZKUYoUDuaF9x/QOnsK5rNn9PRMry9oUwu8Q3rlnUk0eOcsXPdv8ZKJKtIGq4PS8VQnYHp
e2Lhu1nK/Xz6H2dnlwp4/cQ1KgA2TbgEcuLc1m9pxl8m/o14ur53tRMPk7LQrhLBMy0l4FFePuS/
zWiohT3jb7NOEke/mr9S46+CHDK8xHp5rkednQESYhuJjILjwkX54l3ygf7Y6QDp4ga/vltJFoW0
ad7EbuXsmqMWq/J6qELgh0SisrGpf3A9Hlv3kuVi7hZWrkIH9vZnVi5jCUKP9R1+TxAkP+sbDTdE
Emfv8P/hZfaCjTAfXZkSaW7JX6Q0scKnE98JBi0RmXgDYU4F6gEp6E2oOZtObHAEcb6ryjOs03lK
WD28eNLkqjkXTa06cfG0EcuxIKkbiUvad/6UrrtPhxx9/TkFCbFKycsHjxbHmVN8ZRzlusE+XR+I
fe4xbgxY8IdQyN0rnyMQwAA0WnPm5ArnJbnmqQ0X5INvq7hCQ91/YSh6/4bMPosCUsVVQutWCelr
kkqLmzdnuOj4uFjxV7xv1bQj7Q82b4qL5mILGle8in3wuF3sl5vlYAmo9XJ1SXWB/H340piwAjXW
5PgUINKa+AjgJGGKfy7zEUVmNIVl4reeTzUemSnts+D2CZ55rkQ4LI/sqquCwQWQETYL/kC089Km
iG2jbobWu9XaQ0GEg/VuF/F9yMCNSmQ2K4jy87NOCu1UvJ+SenZzLVlOHv42LexMjeW5H9aaq5f5
i1PD4B/koMea9I0jnia/jk21GtCuaMtpjL0KosteEMc0rFKTUFzCbnc00K5Yfz+Kqtjbda9JVR5s
UVY6Z3kzLInsFtokfU6GU3qdwJP35hO3fX4uehsG5+tDjCTQ6JUKv3oER9Gd6Dq5ewN9X8q/oPCi
TpXXQwyE0DGVvwEqJDB7Y5AUaewz0l0NZGOKL3iIXXPnEbKmFSFBPJ7TEt3HyiPYr6bQfLc/C17Q
FlLi6npxFLIaQmZyJyc6zt/0sxLbGT/8iwZUrMdOgLkWzSLSoIuUF6H5A2b1Rkn0L/pB9CpGalST
Nppe01skCAACVM0fypfRL7hxAK6pCW9KlbwZuEDvgYRJM6e+HqeqitXgRcePGZ7O5Yn0iUdjSZ+Q
mnig6jC8YyEWRMjrqHw+8Bteefud11co8FQ40RmV1QEgovIsYLbjdCR0itMSredqRB3zUtddyqFg
Ub0xxtcvPHs401C9efJkZ57Vvyf2CxmbMCFevxh0fBP50+2WD3OKkizwEUBqb6pQ3XDR36XUv/fv
W6geQbRMFfe0b8EZLUdS9mm9P8/3dGnI//yKGfr7+A6VmtKQFG6dOGYdG1NxVHov+KyiQcJ9WoZk
Pw6xtLhqw7cfRpyiTrLQ/Z/kC0JSUk9K2fmZtXbRohNv0WIJDKwBE/GND1FytgJEDh13ZSmNWm9i
YXHKj8QFjd876qxJG6syQASVb5SbLJ2CDeOVGmySxjNLYYYYPz3y2zrijk3Fc3ztpxhcWvikxEDF
7JXThfNcb6DYEzGXojoxi1pXZTJuBuRuuJBMu1+Vys5wS++Eg1a6dRDp5Q1KmlEzx5bDBo3hXVzt
Xvhkmphnu9THdPmCxOyotVtLCbgYiSEVQdQiGdppLC+4tEcwtCPM815O6sQ/3Qq64myCONTBJfsf
19lA+y3jBU15a8aBI+PTbPx51tMR53qciNzL0oPwmQtnJ/64QfxXGEGXtJMRQjo443ZOmA6r2CPm
bpsmNhiQmpkCDs8pV5o0mv0OSsls4qYpXfy7gfS/P0+RVgFjCXrMbhQI9ZpIJLd71K94KSv+C7/Y
yVPkYJ9lLtS5jbz/RPMzOreFiXssvJjv8jbgyA6ma946uD2Zs8AYAIrwSk6NfqOUmGQXIM+crn8L
EP+Bj8UZC5lilnJHyZDe3vIBjrZwnlNqQGaYd+8WpHBlsOdOrRzQitFcaxQn8+5zgz2ljIMk02tM
qCqhOmpLGxwx0havHZ6soHeaVm+kHnhmP6GPhuHGmadgYImINO/JR0v0TmQgHHJukxqDevZFnrpu
67vY0SkJa+1tDRLb/CXkxVHvq4dKWQr+XGUyw2pXR0q5XGH5KX8Wzi5w7fS8FvT2gQevne6x8XfG
ectlSMzsAoer3MSJdMHpGm9pTeX2ni5K0AEZhv8/pdRtx6cmef0Jm6uq7FsVUfW1eeEV7oTo2ZcT
t69LS2eyX+/yFp163aagzH8Yjb3QC74VgmlEaOfe8u9AtZXHvhadx3rRlp//SvV+LivHs3iW2K/t
hJgMLzahs0OBah+28kd4VBHtcqUjMg+QmyG2Kzr7ivh7PmNJMrDNfyFXIALchUmIxKQKRR06NlVE
cjFdyHZ2+Ps6thY4/I+1JJ6fyUkhQwhX4zAB5WG7urdcU/tzICLTV8AXIu2TBaWLh6y2s1wSotXy
2+/6TQ4v2LBmJZ3hzzzM5CRbN2/dF6mslKYe5m21V/a0ZgwJ5Fz+gH8EpZ1v6kimXKSBVKBMH6Xo
v0nIIBU9zUZjxK7yoasXt0tSOQo/M+XHIGTh5hzsH8aHUGizEUtsgalasjOtSTXwn3oSvC52i/i6
eEEh7CLpR4j5lgqLprnFnxxBx5ZUjuximEVxhkCAD4oodAUQRj1VWdNcw+gTg7w1n1+utwqjaSn+
1B41l79+x5PPvOCAV7On3IeOwQpzaqSvrizkwGc6iFzF7Chlql2ljEiS7wg6/Sk/c+TIHUjHK/Gt
S//QkJKTd8J2ojLF9JmIipv7ER+o1PXOru66yfBpjBaAhrAR8ouALhwO+GMzTaBzEHs7CTq4Eyn2
62GL5wpEmww91KkES6qdqLFfwRzSeSkv3e8nsC02js/gj3McdgYvUXtkzV+XOpz6/iUs1YTn0rfA
hMngAGFE01ID9Ib3GpomctlNMzoGjGCrJO/Svpti0Trah3aKoJsDYu5kssddy+w5PHQ5xzDdbAUU
d7wulALr950Um4vILv8b7550aUJjRj+ejYTaKq5Mv0rG9nfI62cV6JIuZmhWRlUBawwZY327/Aa3
zP0EMKn3w0WL65Zq7Xgl556nvfEWd1qBAWQxBdKH9Us1bVqt3KSxendxIwZ7Q3KoR8TFb3WrUbvI
/rv6jBO+qMnKYc37iEYBOWhOaD4fol4ggyk/bEF327MgPOdjvYB4Ra3l1tkSgzMfIZlZnruwRTi8
6bj8zaKWlIDevuiDbyetzuG+l8LeDDHx0HbuwP1ECBe6OOMZ22CL+vf1EIahTL2O/2V6PPmlqFh9
uIEGQZYZhq0ZzUDOW7jI/NRql9eynLtAckIw+WpN07BoT0AXfSZ0DVWr3tg28GUuqW2YreCMNPhj
JWvjbtMCn/E4fsJenvicuYF2jqvhVNOP84sMRoAhoRWkr4gaqjKRFmla/0O8b9kPNvhOmCFK57ib
UVmiDYIa6yczLHQ7rhuk10LyNiPNjYwgWsD2xf1C0se3JJBvsGL2L3e+8vfe8h7lKuPdBh/ViVKS
7Hh8Ozc/c+u+DYYLooSH+w5BeQ8jvSI88iq8eV4wn7EeKw8HfHQBVcdGgD9iW+8226kswMt85Yq2
gPz2LQ1zxWRUjHb1S2YSChN+PntbdcNNwTOfzZ2pvwb9jKNwtLvbOMzProw/0i2xH24TSPLTjkO+
H6dUXU437J3vsrtqOHpmnFcWJbaekXx/5cVW0QA/36YBmJ0NHfxsE+HwsHYvslDpCL6AOVLck8R2
lf/Fup+hJxY4PJijJTYguFvxr0H11xGIzYywqzB/Gu1ZFmwNiMXhCbMoBswdijPxOYgsWL/wmqGd
ystUnuZwBHEIZzPURQ3oW3+L4lueBg1EbH6nSBCjFd01bYu30Ok7dffQpAoCmhXAZFRLC5Ok3Wxi
bVFrQ8DIWy9MATyZ0NWCj0Ug8mDBVERCfM2ghJ0moRn0Eu/dNlr0AycYZq1yjcXwZTotOy81hhW0
03g8XhGVnI6uU6ofvODVtQy/Qxdh3zqIt8lii0aSGVW41tnr+1gJNPh3Bu/piay0YSKiJMF6q1Yf
J3nf6dR9vuqUC5a4D6t//HCzflNaKkHyaM5IHM5+73XBwKoraXsS9jlr8RL2TfjEDmCoOy8EIfzC
jRHAv8S4CttGEjv59aiOSF7u5EBvc7bj5v1dp0iLgv7O1BOjtR20GA4kWZ+kZAau4eRLYCT2wJZq
WIwDoMaSSXzyPKykKWYboS2ruOgW24IlBMS1N7i80R8DB6H3OlBQ3G2+XOHoPyNhahpR/p/J2fpa
gzZ0ZqwTDOefabUNTdaPnGBxbYjdyrj8O2FPD/CzX10bcHMX6kNPN0uzfn9grL/7bWNQLuK34i/z
45qG0BZBBQUEqfZTiF2PwrAvju8ITq4Fqk3FW/SMXJkZ+154ZwgWKZ0Mmxwj7NL1hPzysIuz+cMb
e1XyJl0EWgtfjjgKI9w18GeeaP5/qT51ofuu2F71E3AskC+cf8JHRkzMg2HuEgcPJxwUePEfER1p
Pmbl8UVgnvub+mlRxcHXnEOxEtXUggVaZfL2oewhq/Qn1x1raOeY28CFm4hAuvgN4LrzuN3/Wz84
EdvYmcnYPYiUZ8iS1A0AAZbBLRZkuF+wld9nWDGXozO9DjGh0Q0gZdg1AM+ARGEXftSUJ/PQL3vs
SyuUS09DkbstgTZqN9B+Dp55aGr2OVfXfHZ/GT/4rGmn8e4drtgPf8CWIKg1YQHB2wIqbAmCJ2jv
UuIC3UC+OhXDq1mACP09TRXQfjdPolxJ5ZUhA2Ib0DO4HzbKrCs2fTW11Er7+sQPcqRbuK6Anytm
Wyf6k207KAbxfC7QYq2ga60mONo4mUqDlZbMFk8MNe0v3rJyGa38e99dTOBwxIk7/XOQXKAb9FLd
bqgxeZt12ysIaXC0zgx9dCQiq/zVwRJjTZVHJSzqCnZTC9d2ynf2ZwMATps2AEfOY0skRw+jqzry
Syt5XArudmVB5QXZGldp3zCZTKutwanWGNN9CkLm1b/6XRor3lDXf9pqfBHej3paVZa+KGqtwZT+
R1KZ321AHHANU/AEd/SKuZyD19irqd6cWM6Zgs8rTzCdS8gPz/dl6wgs14zWM64kWP/Z7O+BZ0Ck
Xy1WsxOVQHfKZmmfIgoRzsOx9SD5leC3To04VYmgNqcYFwYtSiABS1+ofM9033gNSsn5sCUGI4zW
mQvTHribZCfNZSa3J4zOSm53LhFL9PDVtVCXkvXbwvKQgrvKQPZqwhgKPnNqXlDIDqPRwTkjfiYm
QK74Aur2vkbJNseb2SbsmHjaeT//MVAvYG7N7ZT4vwHpBjh4KbksCoyzqrSOAIsTeGaFY3mNDQJ+
coIfuM/Dl3gqu6lQKY9TlMM9ODaH7or9R5WXohXMg8XP66rrz7Q+eg/EfRkvUye480R4ZLHAmTZi
xEETmjKKPnwU7hwItKA5d6VhW/+DGFHoz4psBVP7oImk5FUC8pCCdhUS6elDlWP3fnfPdUkOfXlI
vuJVRp75ZS5lxNYgBEtSCLjCqVPjrs4H4Hq59G0b/OBgqY6zt0lgEGE67kGPfHaOD/BFlJwFXMgY
KXM/a+tNYIdoLYUOHH2/vDEJseIvE4Rdk2h0dUphpLA2v90C+dmJ3OhbvU7Kkm3y67az/8KXmArb
If0tiVylRPQ0qmo8ctlyU0fYncAT5fiByKONGiHW835qVk1woFO/GkULuZcSjP3sNNg0RgineZ8j
QAilhaA3Zbw/Ez2GtULPb2LYZBI3TNO64T7An9CloX6Bw1YXymXgNED/GIGNI+qlDMphNeAmJdLM
TuHOTnq6HvaVyeeTSU+2UBQGXYRlQaHEKtjFhmQsdIUtdR3pOlY2WG1360+DNFEoc2aup9/IbbTT
PH6clpr0CmZ4auOmeqqTjhBFJDnjjV5vYA1vQ/JToT3NA+taa06OAYhSrlMfbtEpqcv6f8HB9UpB
42SN9lmveG0/VexVfdOtZ30zfUbLeexy9auJaA0n33rVSo6zneou8P3HHUcHi8oJxkGtgmr8CUqy
VbwZG8P/YShG0vV4ata+Df18GsRxAqC3YZMSMmd9JYOd2IxHh+9ArUCIqwKDfY0KTrm6VFZPD0k9
yAw1WCLsAkXECW67YuJ5xzq11Aq1SFSx4Jb28jvK5Blg2nqaIuQbl0+LV7/S+4werD0EZIBibEcr
vV2576w6f7xHuiToj6uKbB5nlb8J4htdMAgKtjlYRlvUn+Rx0zoRXrUqBqw8+E3ifBXTA6LWHNTA
89HU/+70fACIKMfarYJX4M08Q41Jn9PdYMSBoZyhLFGv0ZSxy2uELGON+n39qIlxbfGck6EVBFaP
MzC8sdDgNE5+7UTOVZxjOv/pJfFY1DO4wdwe9JuRNKQe7CeAgPK6es348hNjZQoyHxw9NPsQ6mVB
ytH8/8g8U3AgDNXzQGLGiZmZe5eYurOj4xnjOd8LQtStoI5mP3+ju7BSBD5Bw10z1XPgGwayRLMh
DsZy99Gz7vypuJSFCGZJEQvnn+YeY+McMpyu+U7E/EPp2CjZ1XPBdsn7+IGqG4BvV6eTUsUAnoXd
3nQEzNhBT4d+mDikm4QjaRyO3gr0Np5aEeZXtTnzQ02A2vQeC0y20TBU+Gmftf9o/q3NDIoO4AQV
pzyHTGzfuI7RNMGRzCvrRrbNftAhkj5/I/FnGd5YRZDE2Fd8UUzM3n2HMZyHQTTudTyVXXezXOwI
wAt1UtX6bMXMTPnbq8M8tSS391dVH133WZgMpiIXaviOajSnJLZyfkaupIOktF02BgdTdJE2Anql
Z16krBYdY5JEaqfAcPnXNVrls90tWHuNAHRgFczNKj6dCipehPwwW6o94epwztTHPV6jPHS1RTw1
oi0TH0PD+SGUPK25TKkZf+dBAYvCAmxnR3toa9fmw8SRfGfxElgtOgyFBYk9NVQqfU7AqvddDbF9
kSztK5h3HqwcOKSg6cKUzpJa+JBugAx8LLPtb7Db65nW4OMm1bEuPpAFGrTwdbxsuz48PeuJmKpR
OAKkao5wqQAgf12W3Mbj77NkYkk6LFjlx1kLzNHigJywYZHjDRJSAeApBge/lLs3ddjQkn+ajzdU
KOt+ZVqrc8G0c7qCDNHxZvd4Ps8XF9OVWMJAhCgXiatpBwqgDFPOcBkBWP/z6rRdP3/DWIZlU0iB
kd0owAyyF+t6bcUzSuKBtWqx5ccfVN5jEwjZ+Z0my1iGWqVgxlG0TUJicWfS5P3o/EtZM2XehU79
p9MKUUTPH9DxTwZ+gtVpv8I/C8aUnj/y/OhN7gKyRcR3KLmXc8FNbH3thEvuclUmx10l6K/9gjDd
aR9FqdvxjmRokycIzwW/aak6qqhHDDpBHS/g4i/dqKkSl0iuvlpu/4cnXzwkFiMrgSWkFaOlLIfr
Ie1+vbTuMQ6JZP6NDgsn0LP82bMhStIixk6YK+GtK9y4ZbxYv0gnEmfqRkzfC1Lek0TpXCbHFB2j
PyKFxG8w/ysvRNMMWXGivXI/+514EQ/HlCZGh++KWyAoeK/efS7cFbfOEgyyX++/xkUirkwC+qDz
zKqxp7bDB3/wR1xtlfHIK8/rn1oKHv7ZFdsu5pM1w1epB/C84BJSfLKMv55kzJ8afM8eKTyrgLMS
5GztKirVkKTTbn/RVXw56yfv49QeGpEUA7W1ILH/dol7ykPm8awz5XUnuNWWEwFdMbeABCln4/en
SjHNCHX8/fzxQbIFpV0RUuxnqliVs1tyB/h5aby4OLL303GVYgW/+zQACQib1tbqtd6dKQmj9FBB
5p1DwUCeh+fGYrgmHmSsQmbtd0O7f9wcoFXz2Gg6u85s7d3K4Sp8XuzhsRwfigclIcdRerxTbda9
4+wRiYW349hlysQ1m4LsoWa39WN6IPpYm2sg2FOROJFq/ic60/57Fr1sGfBdsfJ/s4WUeSmWXK1R
h9jOS0DXzUDEuSD9NFcLDF5PPXiHXAwnfqz75hjvGigDUt24pdrQ4ah7Ppc4NGM5/eBzsdUW6bDJ
ySlCkpB1kmp4OuJ8yQO4mS+z/U9qjxH9RMWLq6lx0lI9yd4w6IF70Oh/cIQjtPLa2qiStcoDfGv2
uIraYfAebAghJF2fZ3fZmUtPaFb8ttIA8OqfPOSy098GLcD0GCf7kxXjmhNg7EqKxkpjcgS/rHHZ
nlURTqSwb5TqFyUVMzBLWFm3H/jKwmZMdeb7dJtWn2mmkuAR6OMBEIUvGHP86y/2mnMhBYTtrwZl
r3uC32ggiUZvrw4nogHcAoGHpkS9poy73EdkT8Q4lowWiGHC00SP5DJbUfVvMUXgsnJivyZ2t/WI
CJo9Qh9Ss6ZB6fstlKAYwNaofPjeMALHz4AsToaJmEc2tFRrZyoM79WnNJm6mOwYRQJ+EoT4656w
w5G3SULCE4EerubS4BhLNI89Y96UO0okc//xY3ukBHgAOmH3Y6dbPjxJQ/9GM3IwMlEuw+5bg/FK
qkPU4Z6sCMlSGdUdaz8hUH87xmkcVdUbigjFzx/jpJAXAeEb7Vy3geobUnOym8NUYgupNrJQGKvY
/smSBART+WiPFZXWL8yZjwRRnAD8N0bpVdHWEoWjhjWICxsU6z5pmrNYRiYih7YHZ0zINBejTen9
onQTZV/Eccxiee7bxlvy+5OHfvYvnfoAauAUxyCIos5JFFcLHOseXW0BFYkWADNIV77nWB6mELZT
AE3tNyvuDK01RUQ5BOMMq31Vs4vktxWhleuxI9Y20VTVO22E3VfXinJLhkK+wlQoQF2KlPCkRQ4m
2p6utlxgYhr8TpTjjk2VCmtcTuCjzDfifaSKelozTUfKcqZDNkdzpQ7Os9vyE5YnjIzYU3pjXuPy
5OSsvyEWiJwMnyLVPmRbTBazeA/sdldtow/Bmtqj5BKvnP49QHGFJBs9Y3QdCQ00uSVWWbF1IbfT
bq+3c4BLSXfhfduoTavYNABAAoZqtjHhmTYTLMSL26fTyjm9Y2x19sJebWNNRnSj4vjCDeO6cwfL
ul1s3NwhiLi2cCqe3Wo+/tPWA4zInlewdK7ldLiuR08BEgTmnX0JXaQwZZtIOrqx8T2Fau7DjMSF
Q3soAZQenEhgUBwe8Dl3o+HGYi0BW6q0pxidUqByklmNyGdSKrHE330Z6o5bG+9n6p5uhhbVJmLD
hrqj6SFJ4Vqb/5xr/LQgdql7VuNcFMGAbCFbdVWBPSGonpAK3DxMBd4gaDpxd9WJl4L9TWbeXu7t
jRZA5ntXEC87GnOiL8wjy04QTI01D5VxEJs6tyOhRKApGiuExdRQWTeHkFqB11FXexrOpEIqDYOf
oEynsKVyAq4lVi08McGgGtIm2laF53gaVi29MEiRCx/Lh3FHOg+8ygFpXb8xZXr80dSHiKHfGvGz
HzqwPvwFZGsUCpkI7X5Y9onpotnhzoqWUyIkpdafXS3OsIp3lMRu3E2yc07AnT7n91XQiJKUY5YG
B+UtiGB0s1JtVblk2VgJa1gB8owonkfY2kxwQ5zVJO4dvJ+0wFHtnUZWVIA72aO4OILYZAu+3JJR
a3h1+6aW0OTcNanCtSa8LEuHxY2uzNacxx1UIhad68uRa70QhVlXyjycCZW9NdX0/izujCrjIN9u
uiZqyH4zXa31KuKQQB7aMder6UTPk6u4f8Fy7VhkwTeAUOZPNq4fVC7+95sJ7D06V26OZ8HZ+enB
hGX2MDEkowgfjLU1jnMUJPfkPqHBr01B3z5KVBriLFVW5Y2HUfFg9OGAW8JtuHhxFwrBU0zGypFM
HBi/IFGa6JQuPuvjoDYwAN1KaLcyiGpWhU413uk6mdJfU5Nb/EVm13N5oUe8k/ortMc5ZXDJjytH
jbkdasYhZj3SBMM+L1GYNKtmE74GOnUxbMvUBoGD4ERPinkbO6BqQ0t5E12idy1C52dxQz73cVmW
LkrRmI+TdVqLDeL/Itd6Euu0ikPLO9/2GYlwxxBnunPcn8dqldJ+hsoeELQbl17lFwTGrRP4IWHC
4R4P5rCoeApBCVhrXGotjGgyYirrH4tL9jwaMvP/i7J4p/ZNRM40JBk+g8chzauHNWpjbZI6SKKC
LIfCUMsjCZ3cMwEGmt9QBgk7rGppC4bIEP8zLWDcx/nHP2xPJofAIqpUM/9draPmOniljr2y6pjy
aAJF/IWLgo+P1AnQ/qnHaSegkX14xjVY6/rXX6/VByjpnzVWv4kZdsj337cfNPjrcAoZdD7/BWiK
Z7kc7NI252yBE1nNs3U/EWOiSGTi9vKYoQx8UdcSaqySidi8qd2f3CSiE105eebq/d7rSR9IxFYs
5o/SnKxenL7VyX5+asX+UmPJcVVpb2zXEoIDM3Qk0mHq0qDRt8QneSq6fmi2iKFnRanMMrKQ4Cnt
dUFtJtDqqMXzcRGv3mGpLrw3JXRpOPqa/MDmHjbuZkjawrvmJ0JClJLvi/2Tc4bCnxFmlHNzPfwC
ry26qejlhYA43K3717Sizv6oqtFu+yjcjDsOjmrLWHLlzs/m4XwkOQsV/IIVMCYRhYu52wXk2wXL
izqrym8OzFRBPSgIcsvdxH2zsN8ZWy7swq/jWqRMECuipgep+Ma0VecM1SmfLXMxcujbjC7DuPcz
MulhvG/+RSjPVxgoPGpCRCrHVuwxzfWBBJxsms1qDzSEYZVgRMHQ77nFtXXMJ3SVR33+Qct9A60q
BMUTy/bd8jwdVxRW3/DONrQuct5VWAaGVzxoq5PtQt+bedY74sXlsoj8ShZoPDitkjd0dI11xx5Z
nhIlaBk8UyTmQ+w74BelkRS4foeZ/byvJh7o1A45bLYjgJfdN42lh6JsRSPghjOUqT3NmsHpvnM8
gP18RrxkhzTl44v9jIlVbCkpEYCXaAuXmf2YGvilGi5GHgaHxPgt7Io98y33uULNZSRpqhsQ3E7d
OLGRnKcSZfj2MjVVssOhTx/qTrZ4qGx47QjSbO2maJRinLOcAPIC3MH9uqXrDChQLTKuH+svAWN6
Y6tmtFZinx2aPKoPu3VYsLR1kCClnfLd88KQbIZfT9AsOxE5V/cFCPVv1HLm1B3OJwgbmQdcE3fA
KpodkZmBcabuOWXZA4nrXkyyVQf+lLxdzItLZ6hvrvHic8F/d0K8NCm7UcawFkbMpMX3TxzQBxZn
wnqw1GvYlDP5+lsb/4KHw592RQ6una/zYWL8kq1er7fyOpUvYAluM9gGSQb/lNTWWoPEhhJ1EtrB
cezFOTozstpR7pnqtjyaXVnxQgyXqlmLrQ/J+9xTvEjr76ygjwJ9b83wqh9zkBjOUIXGec1sz/57
1d1kjQyhLzjubWsyXNbky0p/D1OIPGwc/TwiZDshBNelabT1/SFdfiO1N0iUEmRg4Z54CSFyEGU7
yBbN4SzWsgli9RHQ8wWqoUX6FWgOBF3NVFTiDi0syRe5M7+nJ+vvpRd3UN520/zQ84422caNXiQX
YwKhKVzXg+f27UgYX+Ga1FhTUD4gruOpqwM9GyBFDKkwVrmtlR30nbAjICTnnrXqRSlnJs0tv2tg
ifS2HWWLUJiFNFtrVBCXND928ViRj7xwepc0R+dxQHk7N1TXsrqjvUjIl/9ciCkDK9EUJJFBjgpb
QTUBzLkViFQU9rVOytR8S3+EdvuNqreU2Cc9rcrVTotD0kM58nVGm5IcEFRbc7AK6e3cStxfFpvU
k2QFHo9tKtMk6g5QD+SXWK3GlvA3kLCEwJNzmTkkuw3OrYK95bhmhqmxxM48M9Er0Dk4AsiH2Gj9
bw7Ic2t8ru8l+g+0gf2deDoH8KahoyZ+Ea1aGFrkH7ZpWXAPKjmMimX7ZA+BVRu8M8PIFVNmrZ5n
A/mb7iO2nP8n1ktPsK7BHHLiDe6afL605kETsr3mmhz1BPM7XBzkviOcQlEwEejJ/1qVd7vdnryn
MdZC0M1O0RwOc68IsVbiZN14+ISUtvmEztobNzJYAi/XikNEZl6nXtF36v1S0LDgr0I85I443ath
fDRVHQSzzrD63H0tfp7AEwJOMQYuBE+9SubZ0xZfDIrJgcAUc0AJKbFJ3hnxsnbSYoE3L6xitwhN
suAJiqXxh0fVN06Eh+iDUWYjpXlLN/eAh2VdOtcr/iR0sjFUdu7/76qe0/+8T3Q+sRdehe1TNUWN
oJWElTbTjnCLgQhoBrUcUiTIa2rSvAA2suKxxOP4sjSEMksSaDtkT4+pfj8kkIKKfDdvhdktfn5p
Ix04gjpIw5vGyBGIrZY2dkhNJri72eVLW5gM5hwIngZehwMSUCFJCqgycHXNflJOQa/vioUoHRg+
ftcJTbXJUy2+hgYu8CVCFpxgZipAkc/9Vw8tRdZYy43SAZDvkqccoSL2faPy2eGOi2PfGoeTtzZt
D7MUuHu3xH+zWzcSdf6EB8j/jOcTqx8r2sL4Jbroezp4ENycSswBZOGbP5eKBGt5uuHJeO4B8UQ1
lLDsppr5QkrD4/4zptYso53wDEo07XAz4iiRGY79m97Ypny7yTfqNXfh4S+0PZ8Zc2icbA8UENOl
q6sQ7GDDYpRQfdlnunIbgbRy7AUXHZjiUYaEL0Rd/I50sBuFUYVTx7FA9eT7zV+L7vL+8i5mDoPd
XhFaQpjgduD+ml9hlzwu+9qUZFj65klOS9x0SjYTz2ZYUkqXjwaA5A/93rexd6od5CcYJlJQw33f
I5oM4sHwlUM1kTmjVIphYLk+xzB9rNfF0WgZ844hNSFul9vI7MKnaazr5se1UmESoHMlLNDSDeh6
bXRC1rwf9qRKGttaJscyqs/YiwGFZRw+9S0xZVmvmjQQJACDl/Mjd8gjvd3Hv/35h4MWRbUZsy/9
bJSMPvtPmIWkoIWqMDI4VLaoVxcRLVhHzx+Ne0yHrpNDeiekERcLma7ISulJQUUoApcEvQYJXftP
DjEFRhUA+0BNxYZkknUrlIn3xGayLK+/kG3bHcPsfC10lkzPW7H0S6PD05ypj35LYjQgHUka7Qfn
iz6kdQ0diQ1bMQy7oHb6ltfpT5FQYX2dFqp1uXCILcmoDtVRP1v/gV9oTYp8twQu0SCQKvVXliCo
gIPeZ+JkDWF8yRPniAjdoj9OHVJ+Bs6McyQVBiObBSTZuv+El3uFA3bkmFGm172X+f0ws00l8FtL
ARxA1JdN34YRx87FgkxbMil8NZ5ihK+28kyfIJS8Ki0Pck11niahfu37/UxEuX92zq9DM4+UiDer
ayG6Ur1+IYklrpkmv6Hk42TAzMhNb1IZQIGLaG4sJHM/Hz5oo/ZUjB5RZeu6dGhpNRyISm6stLrx
l8C0WkXhpOtR/dx22QjMmMfDjuqfe71nKwYNh5fKGNk+x8XVsfD14KW8/wwXKM8k8OnU3M0/23W4
eRk8ByrY3UwPErlpCMG3Frmx5GphC5Bh3l9LMt2u4xJclyNwraHzDiSfqi98gyzxkWI3CGavN2d1
QY499pZvIDEc/OClLjAVxy5Rh6mGW18rxpPuze8TueR2KVe7RSIXXVHOXU50OiHN46DVoAWlWeBC
fneJlebGPgNR70rsm/ukFC/WOiAJJOMQNv5sqJHnlhR7KJp9W4qZIrbYbbmj+eefiU1qHhAgdmeT
s5l8ml6RwAtMLz9Yg/tTTQ4qbbM8kjVDJv5K1kfXSohkImnBgnpWy7hi0NFUPj3AOE81qa5hlo5f
Wm4DtSl7vryn44EDAyh9X36nguFui/uFw9lmjU+cvCeV9OkpjSTQU9SBKLqc/RKLy0NgXQY2S3U6
m2qALIZ6LHiFQD8v2Ult49S/w793hOpERPSARzu6A2u69dgsCQKwJQHVAkKo2kaNfUiXaZTdIE7M
g5gJwxfUsWBN2h8Xcrc9KnzsCrVrUm6T15HcYdNIfg+ptm9aemNmFuMSiHNQch/Ay6629lwOziG7
fAwJGS0VEDAP+1+Y6mHN5L51pZJzwLtsqEH4onGo/T8bHtdXdL3Thw9gghMTqfX17MNuoYBtxNbd
5+TMygXVbCtbokZWfxgwieqUYf4zVHM+KA2KovsSDk/iPfaHw9uWSbZukED3u/yRJUNWcKgwn5BA
+8m/5dziTW0khbF63Q653AbM5FW0Xt1dDcx5puZKU1MbLYFxWj/7/VtJrH33k/Qmaj39Dzg7n73+
L0kH8K2qWHLL8bYCbThU0G6B0e44kMYFjjolAB41Gc9rdkB4YUWKCTfLOXDJyJxZZATDEgO7uY+9
TYvJAKhc4NyCxvUDDQHganfrIISqvYpofIKNNf0ZXkD7gGqXmb3hZC6FHvzzsJ9+zsXRlAfUliCz
bCXNJ6LtHEDhbrts+tJIJN6FNB9+kq9guvQ3GUuDiYPwx/BrpU2cyBJHiNmiDF+8VBWMuHAo0Ek6
PvBHePrp1MHt9wKQlJzBOu41tBVg8fPPjF/5VmfCNlgvkxGqeV4vq/q/HKfsPc+ycxHFCLHks4FF
6MvXITiXKQ/oCv3cUJ0/ShviNtg+WRS1A2OEntUnk+LW7AQh0WeTDW7/p+mSASO/YTr0jyJ6QXlw
2+6vjLnEtsGzfSRIk9THSPLShBMn63yY6w5HigK/VyHrtcz2sWC46Aqm5tp4w2O3q/u74QjszQZa
S/5pMkZH8BoVYF1wuOaKVOGO/UVBzOHlvEiSaS9RLzLyvph+8NfVzplDxeMLmHeo6xKUQ0LXCfv+
2yKRj+gqvMnUwQAywtKASb2avm5xizKtsXSoPbAaylCD9c8vkOri1E6yy8pug9L2bgO9GcuXbrFf
gfXWrUBFSiz/BjOCVKINzwcZYHop1/ztUJc2LJzCQBJsuxRG0WtCPDTEoIpuALnykxS8xr07fNFf
umZsKY/n/+nKmAEY1xeU6ZhHT/Iv8MeNAhndZyb9UkZWM2gu/9mxh0N2N/sxrAcWDWZU6Udhw12T
lcQvwn/U1sGigoiIMlGP/IN6nHL9eRwU0GN2ixTmV4hH4ttRTMHL3iFsGb6/GhzvH+VZg3UdLiV9
D/fnGt5KERP1qQhHXsizNxvay7SDEL69qdohGt6pGcjHgSCFmj7Wc7IbBC6md59N8DJvgb9cB5uD
0b/HBrIPZx5/fMQ1Ci8CKh7i9p9Dttx+2uVQclwvKPPodfi7EiX9sxvIJDG8CyKtc38WxmooQWpq
t768HWZL7rRv3tzU9007bGlRUxtn/svuvS7nRuZYH07AKMt4FW8KzpRp7h7Rc3CSEuASpufUbZgI
DepDWS1jTjYk9V78wPW/hMX9bXlXf0NKSTIVDVOpwQ8b/69MkkSeDux1AM4JMoqj6k3NTvUymY7n
BEVyeh2gOlIr29CJT0hmlnsLASPqpkjwTtSHKe4UgsYMSzDx2gKrjx2i2SQDkrUSC6Tl57F+8DgX
C2p08thvT1I3FQUHiJcZ+LMksvJNGKipCVqsF+kftPqAdrVmyi8XtPGvUW2Z3tp3fe1lO9mj+uuD
InkORWN4+/76jx7MsVUkJ4aa4N/cmwvD40XGKiQqapSQVKA60CNygt/AHdD+znNY39lqf2L16XaZ
3NXy57AwfULGY3BkW++wPCUVjiXzSDo+zaauosYxIiVCz0qrDlM1FjmIfkVCgdq04BrXm25g/OkM
X86O5LgS6+BvNNwyCDS4dLnUMOzQUnQsKYMtVymcVBVLzCuLFOCnpZq/+xLt1RDWr3ICVBpgpKrD
0yplq6x/+WTwKOvDTj3xX6pwznKRTII1AFoZc2Y7CeOSKra4RJfLTRBW/22Kt5b2CYmJry22J8Od
2ZE7xtxEcWywz5el4oYsyHMtoDD012sfM1mvyTJgdUOuWhQdcFEe2jL4SiDANCJjYF/7A+6bKFeZ
Rx0J0jzu0u0WvucfkV0yg26wSyRUeGobThLw1ae33HRuvPyKieujzfuiLMSFHR4Qxj7UL8b1vnZw
stKPg+BEt54lpOmN6M6HHHmsYD+Hv5+QSs9y237RhQW9nn38lWmSA+c7+YxUe6J4WRK8JR+1TQYj
6iaBzbWjPssn4kcQYfCYMee2ccaiqZDqU90sdhr8IzCisESUlbrttFQBDXOY0ZweSsLlxdmcHDZ7
jkTCFqd42/+QZU13BLA3V+ip8bbUl7wRUA+Kng8xGTUl9bThyfWBEQ/jz6syIoSb5ps0Zm1O1UCs
6K4nhkRa0J7k5bAp2Y9jx5y9A7/7d5WzQVBVo1fbYiY5/fZQ8d8Imx6eqo/ZcVpo36g39WK2MEx6
t5ppX6C+5YM+Z1e5m4kLyL7748LV0oOQCMtB7JU9URzNRg5dhxpxwhhubl1OHeiCz+cTA1dvkhfX
Yk6d+k/R2/zUiWKumsd10IGmjYmwWC9DSCGEa/wMEYrG/nMc7kaaLgQ0Y2CeeGfscfeAkf4YnwbI
efjrsogGBBLHyE6EZUsWv5uB00NK9HV2lm/+NVaZmmcIYk3rw/GY/zSQRexyN7cBeC1PAQtFLN4N
5m7i6RpDYdTcRj7RTBVRi4WyLABxCvsmkdg06w47yRJloZQIIhLxPcVCuwbLlF/bFW9frh2BXr9J
V2XLn/Zx9hMDJWYVQSti2MfMT2N1cJ9DWa5CdaVx5cFnVYffc7y9T18yelVgqB9ElC9NW+L0rvnk
V/s+ngWM8sofljsMyHt2JfG0bOdFrmNtbZvEG2DE9kp/foMvG0OjEVk91t7nsvusg7W+j4KYLcpA
g3urBxS6GvoSruZLF1DPYEBbOk9yFZCbx+VF+jnbWUkBeq7xD9BrxkRcOy6QTgrNF7Wyezcw2ZPY
FAIf7rBCyL41jRl67he34DecXXKMgzDsugEChPdWym79SCX2NQsVBhtbSyvL+37yv1AqKV2C3+0t
o4mKYZ/ib6Pz/G4Lyt+b+rZWcSn7uhPJncM8pkTPON2gQSln3wP0bp+/XS5YjDlm5tSzMAEFEhdk
6knXmoQofG/lZwAistSMFmFtSJWm6KxI29siQISPVl8t2Rbs4RY340t+cqkfYbl5yruUGsF7Dh5a
i+LktMQgrOvpSEqbrOTPgBAXNHRRC60c45CsCaqPVhEw0YarkOAtHS397kBkLmz0WPqOVOyGijXl
J/TNzO7N+7Hx4Z4Xh73jGFo7yJZHS78BXi9gXE3ltCqL0q+J1oJisyuuDLpZJtBV05hIT6/Cbx/5
xgYYYqs0JoRq/6emIEMGvUbAdF+199tepNy52PdsaTjE9FVZs6Qp5eHBiNXRNzBmbhyBGKNjk3DF
pV0Ab/C8VEqWv4sc5Ps1YoLYyw07QCIfS1SAPYKhioV8X7bQsUXkbbAy9NyrxX8pPHCURPlcXgdu
KOynfgHBNHmv1icZ6XLyAX5b5b0sA+UexaCKqmDExr9VlLwXP0mQ5hZi9OguZ1t5dEPRVR+9QlVz
Q7yJw9hTj84pC7ELJ9/743yH6mL0mPkMb7ik1oYZnXK5Cu70gnXRVetqGg8KAvNKOTYlehjifW9o
8kda6Znid51ZxSUgpJ3Lci5sB8nxtbWaH/LLYI++coSAB+gWW/c7eFZ6dS/bboCdAchLuQt8n/1Y
DriCa3ujOAh/bE5LPZmCO8hyjuNlAolzeZQ1gdF/aZiWmhyF16lC79HlWxfrSNTF5yiRZi2CFmdk
6u6df+QUvc346dnh+I0ODwcym7b443KsTZXvk70uXQxQNq3z3RoJq3ZXOliY6kLSrxdlahfEn5+E
+ia0bL0bkIv/hTmLBFM+pfS2G97jk4fj3Ttgt4Lbdhd8ysjqtRrzKVWnQ82OWNreU+WsdGWjoHaW
+OxP5FH5HZtOGIT5EiEuRilWU74VBlRLP1GDINDp/DIgx3sNzZshtUdynPkp1ON7S6+f6lUINuqa
2SBcokYg8JD3kamiJhV/rJ5c9exAwg6daBr6my1dESnhnqmwiQiyyqqMUfCoxF0HblunSy9eF7RW
459g49KXk+PnLgp3k30st8rTyBiPX2kQBkeMa3akfkAwucLTKAYyse7uj/M7Laje46kPqip0G2R0
rxFjp2EjiPamzd8BrA9sP5JJM98t+2hxba+l8qBfyIsAMIQchj9pcjqVeue/Ot60v/5h6sHPzPhE
RtUPt7xDfN1+3hSlUyNt5oTVVk4MYNdoZW06Bar3U07jkSWKLX9igUbs/LKeBj6QPJXlorCYR8p1
kNfYXVrDo0QRY+5tenCW0ZQlv47a8HhEL+PiNSMrztd1cwnQBlKyGjQ0LMw+50cJq1+0vm9H9SsM
kwymdJa0Nqk8EN23POVwNbDQApC15hYj5KhZA33NLvegjEoZEE1U402iWk08floXLkQ5iefwdQBc
ePxkPHWWvetZTtBMTi/x1UyiEhyUVEF1vzyLgs5Tehhj75agNC2bOK60zNXlAe3PVXO3fm+Nmx1M
Gjn5hGJOC/QaFWfxehTCYgEOYJ55xiQ+KSbmnltnUp1L5TNlpZr82Ozg1ZO5t7uVJy6vaBYVJeAK
G1dgR3pA2yWiiA68FmJ+ViBWFzjbHQ/3dLbkUbdTQ7C3fhnu6ru5PeCNnvpuNnXHcG+OnCBsAb0D
Kgg+I11iju3RjxRSS0mOH9Jf5sIMYWCZc4arEPirAMc0tq7OoVhuvuDfaIA2RuZv+qkp9VhSn0Ia
GGkjFEKn+11dGTNFlpbTFgLrnOYRpVVhr/6H76u7FGUQgx4CyH1wxg+ghqjHipzwq9l1JnlCCpSu
OVLYUsP9V6FGVgbw/NfysiQ3Zl/ml+ezwr38f3cB7FBnZjH07SMqC1ccHSfA0/pO6p9ipUV3qabC
y7AZxAFMHUJC1oGXQvsNTgbksA7904JCL1AFIJf24iGlAxkVQU7GrNCs9Q7Irn79VFUe/1HH5+LB
j2U5pYraTDV1gGofJDYSTXquaFexsq+Abx6CqUdJjeST0RyMmWdOIECMe7U2bZiq5A6DKjX08irm
nxHdTek9wnP0ju0xiUCqffW9A5m3AxHV/b9mYu9sVBuE2D4HcQOH4cJKarNWF1EuxySQqb6YoGdX
Y1xJVm6ziD1kWa7731kt6GZr99Sfpzc6Fo/661zF/WJb6v0flYwmayT4A6Jn0KHjfMeNnjO/Af7c
U0jNW9sZW1wNCivQXsXEATUhF4PyI8QWb+xg/3dHL5S9T6iDoq88tGLwbKkyVRG77QYCGdWQG5B/
4jUxw8glEnEZQyWCFsqPY3K0I7ordxmksz8XCR7xgMHeH0+P/OoOuYoByEv12hxxs3nR+b99gPCd
J9E7ASTPB1Xvvygk9iUjjMONdkUt0sIfNfKnNUVh77lTdIdzbV5ga+nbHwEuijnTazt/G9rwOm3t
wxQYfLYFq6FbQ/KZDqPgW3bAwSJphu8r5CkMZNpEA/yBTfko5nUz5+onuzp4ESugVrDvfXlOJWIg
lnL9dkL1AhsOdnbZIrFA9nVpMLzhbeMFTVmdh7maNo5/lWGYAlYgNw384tp2Rd8fQO2yWiLskwKB
KzhK8tYiTeneE24KsZRBREDATbj6I4L/dmbW04z/uvdQmXGRDgrCyuqncTCbuL3H6agoVr/7pPq1
MK4lwmTyHH3IT40PRPTfqtaaFmOf7qT+bgs2nxEYhP20/ADPvma/sK/joE+zm4VQSjCixBZH4pal
D4nF22LUC5U6SWNDY6PIYIJwl5F8TWTjT67KWKLPsD0D9Now0XbFxkJ8haBsggnG5bdB/lHoo1+5
i89SLui3huTQi6FmAP9KkyT3PH2gabJwYDEY6P/BlL6yuk5nuRk5XU1XhGGP+b79j6RE6OZFd35/
aNYxW8/w0D9MDSf5PaX/qntLq80DUe3/IcbpsDXYwpqquwqKZrKc7FWwUnlR+TvfjDeHVqYx5Y0l
vyKs8KzaMPpNp62V4/Ex2hdQdj6JJREorC+8V9Gf6/HaQ25Mf7wXxicFTgFGf0EjPHjF0v1wDLLB
jrUIVtgEfp1gJfpGHZfxcir0i3jmBq6Jqi+VWV+QivjduBOpyiQpoBzhFL7fUwcycm7cC8yyBhff
f1EkSIuwjAO8jJ4hMU/QtqqW2UA2CVDMg8AErbJrrUAJxLeEb7VerGcsG0aUsisowKpVscvyZUEH
31g07t6WEFdkVUqzPAnW5gIr/B9Uv/L510OUbVVR7pIvL9a+GQhECd4l0L9KzJY6tOTOYYnMzqn7
spAt4ur15WDbDxTtIKmT7YXiGH+5gkC+j9MoMWloLYiheToXedJNU5IK76bMEgQHSN8xWM3kwwXI
KF5Rt53PgPP3W1u/bdfDEG/UK2ANeVtnh8RSDP6nbQEw4kxDEAZy8VMXieZF6NiEwDfEobj9i5qq
33QWsPdI0UGbEyeXu6NVsZXMIei3pkOPaTGJ8m3r5aP1/+oNi26ayAsAJd8RIazQXze7s7plHE1E
QXOvmPHmeNqjFDZvxZT60iBfxt6H0hzbhqf9zRcrmmW0XlVTilkdl4Bdp6mbJo+QaQv3TbQwI7r+
P0tXrpvyobRUcScLpY5c4FLz6dkPgb44Fcq8R0S7bWlEfOIoKRdcmlK1i/hgx70qqfA6ZeYqUM8M
spwp1en+ytZ802jyfxXY4C8Pbuou1C6tSv5xkQ7IU9d0fok3U887QXq0pbkgSFBBiiwFrJ1RYuYy
1Haj2+tAE7xYGXV9TG+1mwF4My51IMQwR3+D1txnLZ4rQ6jNzUP6PnF9WR0Din1OCsgdp4e/Ik2T
O+HnnKaChTE63mDh6KrE5KXayiCfuyZELlIuYHSzj9/7zB7Luun5ryaW4Ia7byY5zclEuqp7abQy
UyuthOUt37NYJv0TnK/QQaV68/KmSNr6NxB+hhHPRhI30hzcEmskz+YSoEaKEYM5khU/pBCAjypV
HTmBPNZ2smzZpcpfu8gTM7Ld2ifo0bwGKhAW+WxNkebnjjZ/o6NhKv8jHHdHBPNTGj+t40evPJHS
rCAFQwMdMhQwvrOzU/60WjQDkf3fxLFV9v6ThZ4xmOU6q5/eKU4ovZEqO0ZDRsPwP8cHuywE26Ei
I5TEFg+jdpJSqjIAu5OR8vWyoPuhNtppQwGEMuV+3PgJc28ezHuQjcStWNEmMbenTZw44AOYQm77
JkDzlVNQzKOxkzwmtd4dd4ihUoDevP9pp1jCMxqCaumWGEvcBtlSJv8tsfn6X5rwNDoaGGslq8p8
RJwoebz1HKiQ1IPe9aUpC6b9Z1bqytvMiYTQZPQBe+eK+sZGZcq9hf7cs7Rtu5pZBH55HadOquKl
1brh13SFfSDUktBCk9QaYMWAdgy3bPqXOE/wMD85Ga5fvn4AyUwta6DRhEwZUYhjvCIWa6i4CiDG
ntFf9C79YOTod/CXw4Q7rrXABK9tws/iqboizIohgwxNvZUfeZqBBsRGEXQ140Crr+LG81TfiBZy
VpNVs7h0mdLMVsJGN9cQHAS2TARln/EqgRYiAE6+mHo1ILvugyGoqy8DfaJRWWWL7G1Rw2KVIRzf
TngI6sWJJBVzopLWpB5fMNW0jKkaHhUEcVnik784vqcl/UA/JoYnwC6qylXeR/Oe3fqSK8ZXCAbZ
aX4NpTllY2TZSxn5SbpVrM5b0PkKPFjPRVYUWrEj399VaI//ESfkocTjXgWqXgq8ZI9tqyhGHDmv
Q7dhHcekthnd/bOSZT7MZiiHEG79CtYA2dumg1fq9ya3J3VZ650B1VHhXmWPxeNA3IHei+0JWEdt
24miQmR2UIjKIaxBrC/l2CmZdoFKnMUY+bGUZUgC6pTd5qKPaLuh/55snMe0mNHaO28LZ1Zp+u8k
L3PhoWJ8JlYld2xs+sxAUyMCnloz0VVrg8lk4C4FMD7gwa7QVpudJqYwPo+My8xNvwjdpnaK1kcM
wv3V/iqjycu93EX+xfHMJsG8df2+FxDKBOi5/0ZNFB6NDL4fxq36AiKW4JAG6mA6Je/9Th1YZn2L
ygaAOIEGLEQsg1enlEIy6QC5/BYLpbHQSEjmNXajO7WQFwIeW/U9vDluo9BpJhQd/PIVwS1wIwkP
gAm74uyt2YCuEkwD0iDKeR4iUPRN8toiBZ157aomMwSrttjo4V3j45OTqE7bRyMztESmOTr3R6Le
p1rVNjEzyzHEBq5zAqgtuOmn8EwxV7U46p+NxC158EtBJJ47+xsyw3j+8i6ZbsNf8FermNUSmyw2
8ZtDnnqk9sfNKisXPUzRP7oredpKzo4riCeLagxQ6TirNH2Tm6/0aj0OrxZRxVeUtF8Hk0glzcOR
0vXZC59vQok1z7bOxLhO9Xcm24UdupeaA5YuznP0i14mxqztJp4lIldFA9P3iZePji9kKa8whcq9
p1ysJqw8NFY8Zce+MooQVrezBF30pnhHnGHSEypROQ64xyobcST037+AGdLpSkQGjTzZN6qP8vD0
7+/ht3HZ5RRYcwp/oENu6PuxK7zigSCWwQtS3H+T4Ay3Cc4e7swFmMfWl/TUv03vefmSWeOBxGtW
2ndDp/Dq8F3qsbbQsMjQkY7LCj+KX3W4ve/aKpPJ8ZFuugLTsLmWUgT6Ts29sdLHJXaECC9weCzM
BYnGQ504Xuei8Q6vHMceqlWtghXqCKZE4jIggMCPQZ3SPGNakWDsbUwOzy5eK5h7A0ktUjHXkPG9
WitC9x7GkLqb2dgRdTBMx97F2UojZyx2rebnI/XIF/aEIk/zL1d8HbVKJjiDhJcQ31nweGgOnl8j
dq2zIZG5WL1dnRG8x86k2fvS9dgULlKPZUPV51ic8n5TZzKE5erZzGl71qzYtGp+vDJVKhNgfPJ6
CU2W0G/NnGlILD6/BHJb7BGs+2FA0GJxSXnbrY0L3B55+H4XYevgzCXgFunfmAWS41hZ2s9TsGxj
cmyP2tJxnGq/1Oo4cLwMbMBmduZ4pA+GRsqIYKzsDP40jyJSedB3KfRTrsSRO9gXjZkZxzuQenrY
rDi/otY9xRGgqT5QIWFSLRunz2/q6dX+99KnSinh9QW/Du9A7c3EwB4Zrg5nDSq0XOX5LsvB4mi/
2Js6idSwxjmxklzpkTuyuz6Rb9i3yNndGKMWIhOT/YgGfQMnabGAnHwJsxrFD2Xy4TWEUSwTkodS
VlHGa1vFxMOglAxkADFvOnMFkU+ioriRFTXqSlduIIO9rOyuhQWZ/hlRe3gpN0KLPOLU6NoeY+kQ
ZMCko5qyby/vsXhO3l31PRkfRy4nzUkRWOOiE9uoykUHvj119cyhyyKsH96x0NHnRSwBG3xS374L
N4Z3EKrGZdc2zeX0WAZZnXmrTq9g2rAlHGIz3DI7RgmSppV0G12r5TPYArSDznDUlpPlBIFNp4vM
RI3JT/FqbobQxTPi+88WF9TBDEGwfko28JaVgqdBGnGQSKbON1QW8aH/dEgrLfJqnvKDkqrkh91X
qa1bOag1bEgy1c/D/hSiEwaT2vNv/puiXSEavbPAyeWWA4hNWQko7kOw+rKXi/xigsrPEl1YJr/U
irWFfJLwIaWrQPkc4uuXei7+mF6n/8ku6gz7DlcplJNgsCr7idat3+O5ZhS1YZjhScRIp6fKNoWz
gRi9WNGDfDH14BLnvi6xILLpu6VQTbIuORvKrsCxnm+TAUw/fcMfdR8SSq1ytKxaCR/5ZgcUxdKN
L0UPvzHRZeyuoKrYweYFUlORh3LEghiFm1ZF196Yztj1ECSrolBj9JrFa0ngL+FDOIBF9M6yACi8
lItNwer2HwFqN5L7OYR9tsHp1eORQMvMBuxcoj5310JM7zNs83HBCPW5tSNl4tRm0CwnDP4NZYRI
FElLAskLaHUGOKhxpaQPBEms5hcBXvEltq8kCAN0Fd30ZTq7QzIKiV6bSZTRyj4vRXp1gktKKsyu
37C5k0btNOYRPcXs8HzzM2lj0NckaNNH1Q0ZZAKKxN0pFi7oQ9LKTPZaCmg36m7Os64Xc+0gJ+20
yleRZKeKmdUXmNlRZTPOO8pyAXOZFXc6ntHOASXPlY6BHaaQ3cd0Q/TgiW+S8tC6sc8PbyAQLv3D
/bbC8fjUPPkH/2jvWjgPo4k4iLSWLL6oKZ7YFPVAkpSb8l78w78N6SKS4QyhQw4bxNB5CYixures
9DNb0YTKNTpKBCvObaGQ2xVcT+9d8Q1LE+6ixlxyYt0xj3FTMbTzPp91OJ8wxyiCsldq8yj7H97A
zrd8CPlhqIjhKAe3QEIsHRKQjVwvFhDiGU2PCr3md/wpdEmZJ0eR8X1QtT7+1nPQSWeioGtkQ7+3
o2FUDuxluduN0g1tcEw5Bt0Jq/zajww13tS5rG5luyERU6eMU8cK+13iQzA0b1dJZknedfhKp3HU
/cg7EKnMZvKAHKVMLICVEfWYjO8gLywjxQHtq4440WYrJmxVLHE/sXR5yuwnmZu6isSBsIbbXos+
z51/dE4mEoOC4+LswMuY3xz+pZZ3pnRytCbt9XpZkYzJ3AXrHtiCqe4pC2UkuhvWzycYgAxKdjHV
fu+HgnBfJZha1iUslfZQfAdmzkEzHm4oXMK0BKpXHFVZhRHCW7I5E3eeUervEm98M0mncuIP3kY/
UE3o6FozJMBChZiOHjrN3vTjNX20PZGyFYzyRqVoKRza1YCCiKOR/fmulxXMCUy4AvGLS4WHQAC/
yFwb6/KR63CGw34tCWtYjhTpyf8IhhcgDuZ4Zlk6r17EkIOff2GD4EeCrZ9gIGPbBFUcFeS2lsFS
+kBfuGRCwF91MVf/O01OQO9zK1s6OrgAAHIysswfyF7gMThgBDrJYP4PXfi43q2MuJk8WqcSVE5x
grSAANxc5TXunhrqD9UpGQGcjhGWMSueYIpfvCGaUGSNEhdE2q8ddZoDeooNuAlV/40a+/b5OKqy
kd9O6wvRTbEl678Aze8hzDflLhvhi/piNE77DJqZm+VZm7TdmSaDPdwuL5Q4MbPT31HiOhPmg5q9
b6KXBAbdnVdSGp7VNOpvcderW64BybhinSWtqtaVKmN3IxJIg+BsWAmde9LrqBJlfKFm0bQLVIBY
YuK+MSN+RcqJnHMdVU6Ht0we3NPwtXwbZsDGMF8catocQJ5hMV5ZtyDpPPbSyHb2zZuW6NdtuxvZ
30QXDvODhTcgiJmY1KmhkSj7znpTFZ8G1MX57wnXfr39WCOl/FMK0eTAdTSpqXOXtz/icFfseBLF
fbsA/UdZoTr9f6BJ1Z3RCoaVjJ6fUcqgiNw3Yk/l3kELyq+Gu8P0HtiHrT3pWwQE2EQ5QbPulxEg
unbDdGO+mmYoVh+4/TFrmiBLiTL/5IzhSoMZYCk6wn+I4PeDe/QcEPeyVfzrwWlZ9BudYCkYAXv9
pGS5j160d48+1WLXu87k7cUvHmWmB3WpQqB6lA1jgngRTzERr80CkXmdff9P+r8A9Dk9trMC1yqO
GMX59FlRAT3FOKrE4+ZLNNf94445GVyrd2+lEWDoykRg/G/bsO9ioZT6HTbs7qwxM+pkxd3wAD6S
bF7blZrMxAdkM5SvxMX0PdiQUVqOsULAoq/TNn9eqwdgBa8WL2vmJDmCm9nEf40RMAf6myxC7xJO
2NOl0ldvR40UVXXMkuX/RO8BS6fomQH5b1uSd1FnoDuzLlLMgdN2VzVWSpgCp8KN87HUq7FYahAI
5+/nw/Zfhz3RQ3sNY/VOQKt4qsb+kbSN3xbaB7uQQk8MuXjjVp2mD4ysQFFdCSeY2lu9X++r80S+
nhIdC9EcNG4C7R40F5Rwgc/YziBCoIjdCQmwPhc9aYQnIyR3mzjBjqyB34QCRfgV0IiV0yTWlOZk
PIRz43uP2cCL07O5azntTy5ZPThkexBa8n1zVIuCVxO6bKP8BKTsuQbN5h/ywSDYi1zEbSSsAMtu
oQint6Se9gsbR1wnrcix/ZiBDyoAc3K0/WZEeTkiqrltjGnhVzTV6ciWr1EbFt5ar3nNCQNgmMHH
qeRpEOWVUKAVHwG6Mu6fhEk2CeKXOsVsccgUklP3N1ME27vQO2Pt8IXD/6+1IvOlvDTG7vfRTRk3
IGJVtRPaKMpk401o8epqFkUHmVIiLIJPWDg5Xl+6BPDMbU/9f4hVbPib4KhDdMPsLU+Lqt83gcrY
xjtI0mcFbrcZ2Dbp12Ezsxv3kgpUFSlqJ4UPu2wk+8hM5TM75vPMM7uo/fuX18P/RjQp6j3PcDTk
L7/yNUkW+bXjZtMGJRXSkIPj4FosZ6Kvp7G1Jmfz6Dt7T5J7zqnzcWb4EeUvsjpGrZMEhl6oQGdX
2MfDVc93+wDJESMp5k3bdsfvPXK0KgdsC/XzsAEp0ZYo1vdeVWWkn/bQC0Izz3L6l1yZD4v8ZIkX
3Bzk1afHdFrum7iXmKETeqS3bkU9cluBtVeiCvH7qM/H9AMP3Y8R26OBPfzVqR8HeX+C4oaFqPly
ScJxwsjqbX+04eDHvTqFMEe/zigGyjEwYWl3bfT5oS3yK1Fi562WeCOwzLyhyTczlCJmQPr3fgFs
hQzX2Y/jBk/8YWOJRmV0OWXdtU31d1e8svsb/woFXIKvhxjemaFRM8g7QUqBY1Q067ELik+37cWN
BUu/n4DZmSWxOXYj3+RUnI7zOwtSiL/Par/2tWHkrcU4b8srRhx+ZZXJrbu599KRiCOKy9INiyJR
/PpqUrphipE0sVnTsHuJ5gp9N4s53snBwvwsp10Ka3vCwOBAionA5UG7zkaqCY4tCKa2IbrzIx5o
OGb9kRJ+Ju/pVqKJ8JcoFt/P9kAx21aHufk2dXqGprb2vVpkTZNFCaRIXnqXUtRPqCdsRQGLXgkQ
5Z1sS7ljR5up0LvZMXDXW4o58ncwkJ28t6P9vEJtwt1vouXuJEd8dCoOm+1hroOkHSZIMCSPWI20
+s48IiniT2iFu/sEoc56EOabWk+a0VtHo765WiPZ4nGWg00QHtJyq3g7h/ATHE4sLi9h6njdmsme
HS2Nka9RrYQT8u78OrvCBH4ywj8QYEQihy0qGMjtQULeb+f49W17sA5jfFl9G3ZTkYTpQDm/G3ih
OZDTTz+YkLVOwzOZDkZBRo3KD3Cf4kGWB8/w/OYUa9C6y7QyxqfrFHVQruesRx9ypwsAmODlkpHk
RRoxqDn4KZ09KbgVAWpI151Ke/SkOEnY6phlDZuz9GHiOZA7Md6A8P8dq4lrzEtT5jR1fR/BTz34
YX3CfisCowtEGM1tEvigb2/La1iOwjMjx4YDN17w6RWXTshTV9Rtw3Y4lQUjiYVNrBt5Ibwyw6A2
gMjOl2j2WtoL69TbdKzQgY2eI+8LjEUQRJj8/AFS5702HtBAqDx3Mm4ExWb4phHksfSpKYhiYNto
HH/j6dYWN5Z7wPN2k331QF/83rW2QGyRlvubxVdm9XCo9WBa+RP7P/KJCZS7u2W4zcLai2JeksBK
mbEYZ4WKmcPHvttP0OLexysg1SUGrxxx+s6TNevC9H0CsxuzQPID4vCWr1qKD9EzslABya3qjkto
SNVrmvqS2K5ZBAFWhgD0+ZCY3xqtfIzzCNuWhkViWYh824PvHSBuWfdj41zdcLAo6luIxPtRp0MA
GDt9NLXYuvVWmMMjGVxWFwmPjubrifuRS6aeWG7M+QWZdL3GI9/jF7Eztp+puqWcOxkwAlUFnVqv
Qrc4AgPiYHRcA8JtKzGZUu4dM3nAVfBNddRCihXL2zt1qwacfe9WsKluYXFioIp2LXa66uWTmTx4
GlTsWND4q7YutNplxmK0FaxulLHZTTDMCxWgdII2SyDnXJ4imFafAB8yfhMu4OEQYdu1w33ib5JZ
ED76SHfH9yi1PDgOP8bc3Y4n3Q2XscF9S5G6L7s6PQcFx++UKnlRTXz1y7r1dbGFJ1Nto+z2GHuw
iPfjDrVQXa4fgisMTP+1VBzFxCace3Hy/hXL7CDgghq4fa57AKyJbWrkXaNesR0qga5C/Iehzdsb
wG11cLgopDRxjowuNht4+0KcFVHe7lrTEt3YtrMjkj9NItj9TMjOhZgK0o8M13MniQGuJh3TkmLg
m97xiSPtlM3SkVevwFWKnPIWqkXXHriamAeJdNxyDNENh1WswRBfDkBCkkCgXsqSoBvytF3UbLBW
sFUOluGnXOM3WmO8Ts9/Zlz7gyyL35JFUwd6M2R4cfbMn0mNa/KZlVvK+Akpb2j7eq3wXkoagnY+
XJ5kQPuB7MuLWg8PPucmQgOfXgIGaOduKmAfl1Er42bNz+mpfeLSswf94adnhPZX+LkgkSjXjQMh
aUUQPUlnR+Q+Xcu4s1D+do/rEiH4BcwGM5ZOhlUrbdAe0UgCbVjE8wRK1ac9ZtzVNvSXlwFSTUEl
nta/jabPCiH2sZ3qn+ADve3NyVl4yEY8hIahdMGXkakGcEkw4Hw8vlECfizMvZHnVcuE4b4NJUZY
F3kmZ7KnYskRgNGEBhusVfCoTcW8vfNBsFLYQ6Z6j0ggbiDAvIcdUWnjizGD5LBce5v0objuwFhr
HwzPRg4L62UFkZAiRuunafBXdF/MK5WgM8MC24CbXvZSP3Z98yx4gsaMFDev0fGm2c0Tp/UWYoAv
VoT4ye9BDWv5YlkvA+epVYWcsesdZRTYEugPBwNYS3oVLEhpdQz63UF8hccAfclORgKrOlfh567r
UTc6cGIC2PpGhRLk6fAlXDoB8Qs8HzYiJ+HBteyU5zcdFRFCYOxtioSNVVaC3nHjaaDQ9Uo4JYQQ
U4//aHvImb3L3n4vNjoOOrS0QNRxtLW2bh5DgYvFDJVH3J/1GmVBA0gFo+lyeCPO+w6qTQ+27fks
hK+9ie2RXymXVXbT2ZBenI9EBjuvEWk0HtmLpiUH8KjHjYoO559Levt6vHJ04XMxWm2OXcBFN9qq
RQTuaQiRgwV9BHlRoiA0R/xH3A7kW8JpemeDqDblUeXk/gJJg+cljWjN9dpaURlRRmw2jQsBKTwa
yUZHrXk1xUk9vUH7nLVTSNDo990gTijcgI8xLNHSRQnWufkGx+hmoTGk6IgAq6S89i+73FWun1pY
ZuX50TNgZdav2OJr4yLYpz7U79wPOp5Ix4atKrRatj8DIiOK0T1jPDuSSJSo2I/ZN7cWsvFvmlUv
Z/zb2UXT7I+cNdnEJuVlud9nDNgXMl3OLLXTi8e3GOEJF3QE7nrx3RN23q0ala5A2wnwgaVdD/4H
rJmsY/OZfLueg5qBVDhDYzXnNlvV3ZPQ0I9/1j20zpmi89gmNHByVMIdQBxez5s/pOH44AEeWgkK
YFZuJfjP/KNh+8ypI6KDEWbJY7rKUPcx7wMN3lY7ZAK8WKbPyZ3vh8NsHc5WfDlcaIkI5ANDhJmz
7rvG5MTn7SRoS+VHT0ZqLBr6zsIbRMLw9tb0ZaWPtUj/0zIChZvsuCzO5Y05UQ11fdg9Xpz/t3En
TtURUFSjryL6KLPYAIaxb/6sy7NE/Us7ADFIRmJMwJ2a3rNMzRFqmCDKzYW7Gh7T77dR+7fQwJug
aJliXTiVY1HWXtZlhaeV8XSxpoPEOFtUY3xYz9ak5RNR7mng4gGr4pqEDf+iRASaa6mz8FQpVX4z
h8fduB9m/ZjZCXfUpGeHBZWJrhzGWM3t/RWAvMeMF2qZO0p+iaovbbg+akg8hAAa8M99fH7OLqu+
AZqL2HB7DmmJm6F5cKMttZ2Atej932vGL28s1IXPG1HBBGr9yOoOJMWbS7WpcdDVKcWSdJxnfGe8
RzAxL2P4Sb1kj+LG3bluMt4ICkQps6u/6KONCcBD1nrschBMpObLHZNXgKTj416pmg9HAzerQFOt
QUXcNpYxJJ9wsMr9O34SDljxvVJTOhjvphO2tPyI3noMy6xqPmG8jyV7pZ8xQzBzQd+VxLqgfgax
a7tCs4kWYHz9hxaNPYKFYj3Ffe2jXlYLBFhcNfa2b/GWlgFw+dzK/a1CsGaq6S2OU3NL1nup3A6U
QH7eyYVbZGFuo+1zRdhG2LE20M5488/wjojg7hHd1LHyFmFNxOad0j7QJsevTZ1XgnIGT7ct6lgV
GHH+L7C50rOIqLTcL8dtqHydN79VERHYKB39SMa8bL+KQQ17IUDyrpNO0EATp9AsmBUnEo7gla+C
Edqdcm4AXc+FzxEDPRQ9KMcGo0PjECV/Ofx+vVTEUew1j6hrXF5/6uWF+fFa7TsVn0dreSo+49LC
Lse+QopwAyl4aE4D7+brV3XN4vV5X8u93/0oswMQ83nPcC9wokt+S2hKBW60OL/MrNWksCdxmFae
+kQinbIKW5nL5oK9EPjkMT2WeQQxHZhHfgZ3VEqszFb5xf5H8Usnh53K5kdszze5LkU8zpddxas2
4gi0nd8PUSkWIaB3l2Vx+gucLXNMFdzCnuBZddYY5P9JEKJyRnAVLZbwbDXmGoFOG0HOr7a46yZz
JKF+gFXXI4hv2buLfEZKLKjEpciKAthxpuXNUxXXMP6aYC99aPigaMIfgT3RNW4Lm0Zd4KdQfH9l
rbPf1LBgONcYDOpCVvdTQYRRNIxNw+tihKYRHFlYihaRBQb2236fD1dsVpQ5G2dxK9sDAEpVTbae
QC4vzSxX0yfLEB15PKmVMCYwhRyFgVnGMylgBotKuqTVdCRsyY9IzH7ly9QwRz2ayO38EG/aFkHb
8o3t9698agabFWmbyeclHr8XqL2QuB/Yq5yIXjvfsNrdWBprvVBg5nx77iEcq4TjAG+4lyUr2HsY
+h1fXqwdsz/3u40zPrPv0pP2llfjmsfXNryO0LCFf1Ungb+ntUUmm5afl0Ndg+C8kUHtOUEVFheD
x4kTPUYeqRoJTXnamH8PmZwSWOtMrDZyn9bdS7bG84WdNrr0/nhjlHJ4LTlUwn5JQRhRZcvp4klq
P2zjh7o9iF3TmRG+W8Tb7sux+iTW1ZayBJVbb4VYmJyWMhDW8mu6QdDPQ1AymOUSgjHkpNm3XHa7
pgT5rXAbTpnuNwTXJhnaK7C5En5rq3n56slEm5imdPqvhOu1ziiKfB1gLH+sirAHMVwZaVD3U8ny
7W0QdLocSS7Sa1sw0pr7eJ60yl4Il06k8QlUTu5TktBlCEjbkXBbQ4mcTQ4eF8tI6F3+jRh+D8uH
f0Ezk7DVryrZgi47jFhhzhcfNZ5tughcBC2K4DVRtXs3x7kMIqCOEWyBiw2hNb/ol6QS4On/AJiT
nVivHsGoXvbK0nSJIE0oGCRqk+JXjKrg+Pio65JWDBN/N8lqUnVZZf84Wv2BobDEnyBC+S7dZHc+
m77VPtkuWVlexwFV0evyJXZa9x4CZvsmgHaVGvW2GD6BrOfxAiou/C8LwPTFgaXw6tc2Sqg7N7/c
k4psuNt8J5kjgQ9ERA2IehcbTlN1NaJbvN0tHBxfawf62GjrA9f1XNU54WBt3wFN0oaA4LluzMG9
Mkw22Z4eVCHXFtvAAHlxC/1sPltPfuzmmFn2yGBxidHsN6mLqGau2Ptya0HyHgt0lrlCx+2BqqVK
TW1PYVnp8h/qoL9vubAtyb+U3chdKoyu8hEsRrfKG6/gsn/jcEVigQX6Tf98NY3COM0Mi5XsOrlb
9xfyPpJHKe9x2ZPYfUSJOBrkD0gtxQTUwi4aaNRnSOQEW5O/64mt/iQtzq8pt/a5zAvfaXqX9lmU
B+cc+FQz4MXLUM4sYbYpkztvA49VAlmMlbcbBctWlcIbJvvDnoz7AzDizYoaE/nA/+Zm3BzZ+6v4
Z+2mUa1Ww6xM26aaC5Z2dLGjwAfbD2LNag8hrXfSzqMwpbQUaCvPQJuKyyYkxS5ZqlPMvzFe1INt
e0fuUixZBf1mrel+jowgnCT1/PFqB6monDFhhU7UDPm4cgyLoJYkR0WDLXFIRZzDmTu5kOW9nVYa
9k7CcqfJt5e0rsJ9/pPZHAMB41z2efE2mLxLzgTK0KM3BVTzs3bNjU+2cBzVT5HC78RX43eOHyjr
jBjg/yhxWEMwRQu43cdJSAGcsjebOB2q4GRc+rhHTM77Xo5XjhEjvFMKDRWhFEqv4xdmQMFel+E1
Vl3oEfSX8N7ay+twBV5bvX6OV3PilOR9qDI5SBH0tioLo4sqNEXPA01MjnbbMI22JNG5GSLQZx9Z
Utr1dDUJvrfCgMat0Jqfh6P+Zl1zKvotrma8smKz/VI/eIj+Amv1JATf3jbvqKdHLre1xWydkzRv
SoJ+lO670vn5pnDnXAQS27p2rxLNlopjUNlW/8/CUu8ysW41tRCjyg9UFtvNmEhJrgkUu5t8G4Y5
NPox+nWd+JpIBbK3XGE1oC5iLmEJxyKXH/YYBfqlTE7pEZb5hAOcS2qT+B2pddrlJo9bY+kSXoOX
lsjdRNo+gurMYBxEJLArcixSSWg+NMzmwfAPkjJ599XhG6KE2Z3r7yjFBUxVH/0ksdGvQKYYUsy0
y3ly4lTup1WWiTcVHgmCpJFR+CHYwsixpHXxgqzWPIm8PIKzzvUQ2iFyKZjAwp1nJV9y/JNAzLM2
6rsN8c5bTQmuAzCMTcrJn3H6zwfCfx4gLty1PeySWK+lC8166Z8rwtgg6Enh1BUOhfRB+br0gE17
5GC9wPcfJOFAaDghATspgPCfkx/Cf1LOhaYhasdvF59K10Tg5AtHG5Q1VrZdhZyuT8Iuqd3btJ/s
XWzUaNLiuPs+jJK6+B8J4g9AFrzJ8dcJQFeyvCVxgxFmzlWHAG/ylkDDp9z4kNSKXgIzHw3/KkHp
H/yB30XUqAolXq8gBTUJHxOfodhwx/N6l8YtMYFzU72dGAw8nyDBOivpOd5l6C8GwrAlL/RxR06R
7mu4HVeBSnuM2e9JOYsw3eMRc59OChHkyV3d7Eje2P8yzyMbus83r/DhzhqP/g7KS9oDBxsE9T3x
uIsVccXTAcd+dtDPahfr7a/1aeEimERHgIld3P4UOT4ldrWVyLrJ7Q4TiLOpqVMzoLN3zdmigqZt
sCxThKpV56Ajcw8fDZoRw52xPMbeicr/h1K6XBdV93OcdcbHjxKfFtS42XvuTnd2ksUFRDP4yw8v
3FoV/EXemdAA10qKJzPJYFLGZAFZQTkSy1VC4ilVnTcIOxe/Sh4qylmqvt3JMbjGvF5UsiundS05
tsyXedpKaTAAFQrMeIuEERGw05DgzOzhz+bCv2yFuAnflLRf4mvnKuErFYC5NhrOxwQUkskquQ/G
BB5D2XkPSl53p9eIcMHxawql6R6yGKUotuNiLqdvV5oJ/284JFTjE3Qerb03+TrTFcfZUyTnxydx
RbJwTw8BvP0YjifeUT7sQCMHpNILWWT+VVgjlyz1oi/GsLdT3bRxl87FPYZa/e8topGZ+NhHFcQd
xaM6zxl+J4qlyd9i/J+9/h2Vl9WdnQMOI0GTUgaFaVjEZkE2P2RGe/HApuPvXWtDcfgJBaui8WLw
CMBWu+rKRAxH/lcfQd3BwBTw+Qx/Ch4W+A10Ic5PU12r1kgxJHdbD2LXJI0+fFTX+cp/S6i91ls1
OlJZ0VrnwheuwdPFma1GAMS+MBhqiVZsB9U1zpSNhur3ymAOuFtEAo400i8AfsFo+UjKadRIlZBj
k1TLIyfarA5rfS6kVEGM4ArFUDCoO4+xxBy19s1jVgUyRTjEsB6hYvMPmqWrnaPR7teAp0DW+nB1
cWEcoI4CmMJk3O73FFvXLXBVseBskx/lH/oj9Isfs3HKwqvmnPK7nkwlCEwPqv9kYGOGQ32GRUzI
9DOenyJI7eS4rwFvPMz5kE/HccFkaARDmFiCeAoWcouFdxMu2xLTcutkpB96C5C8Wdmz12pE67dD
3eWbKNZT7YZmoGXsfRZGyh7K1GCgMJ0OJtGLVwAcrleaWy/4sbPPNEYhSP4OOREWvv7VznloUwN4
OoZwOwZKPbtwBT1FlLhPEAkbpipJGEk/qACoZnmgWWWmhFE6CmjjWyGLS0GmDwOMx5+hZcn2C0zS
JADVtwouS9rnUqBecQlynfgqFqDgW/g2EkfjQjkxslwKVhtlGHfoeXfWzy7V7HMv3nTAgtIUzzW3
ULIZsRekuhGRx1f2ii6iFKSgAlVOjYegDg8sNLn0ALaIY09v8cwJ3ZcYMHC4Jc4yo4+FdTDaOyer
QV2gCyQNIX49c+Pc5bSxcvwkdF7FpOAPFrz2p0o/pHB+3MHup7P+31UNuRkUu1OO/QpVRaRFX5Ya
/YSI8yJdHwZwHo1dczmTm9tVVwXFgSuBPXFiOmC/pINNs6D2lz/oRIg/p0vIXDYUQjYwsyCFBBur
YZujwYfLgcWtCpgFyiDc4yxYyqOZnkI/tLn5djmEUua/s/MXnd2iXK9cAmruZ5Da3mVTX1ZGHrqg
xC71K3/LhYXaK/rfYjbC/dG9hDDvChjhNZ2wXjCuZ9Bibd+gjykR/okAv6wrY3LLiYA2b+TNuX6c
JiD64i1fheBWyKXU9Mq8xMq5kThuUt2OoxjtZrU0AB85z3BjnCQ/wIf990Ouuf08MtDK5zfbZN8Q
uW6fLzc04/mxjQrzMo41DE4NWoveWlfuqvXpgMnAoN977WhgKG0TWStl+CZ3BhlgeYVyh6FwWx18
NbCg5J1y3Or3BnHHB6GT/kMMeX0aa4koKtC7o/NyDE8KGNhfhfKDXeKhgU6anqD3cx9cV0hCuumI
D3ooU/gVy1pculNXbXG5XfHlVrtpJFjQiJ+mi5svEy/rvyYLsONMyNetw+yyyQVT+zEbzhIk4caA
VoB35mgoiZQ1S47o5OzcH7LlhJGWFJzI96PMD8d+Yry9qyWVVrNDslP9rlpMw7Ctm9sDydpjNWpL
yTSfNFNinuKQ2UZNmXxsxOQDhEpfQ6AF+j4PvMfFWPW07X1DvzNkMQx4y9qt/+4rfD0gQrIseMHF
6EThZ3VkA42Zg/9vhghNdQc4/YOJ/e3KKGCDQyid0CyPGVe+p1S++CUtO6Wa8Qh5JX2n6KB58wXM
hOVpxUl/hW0hn6QKQx9JlNXq23U5Dubur+52ig/nYz5xp2J4ZBrOAVHsWliOVG5MbNxR1KRP9kUK
430PZDCs0JahCUUsNSW51q172orJdg+gBqXCNM/+zHE1XtLCkUnHcSdpO4AxSLFzR+KA4fw9eRul
C2anq52kTdUdl5NQTVOnHtPO426nDD48gkY4kxoboZZfU7bxvUM+TTbPUXK/6v7Dmc50svNrlfkg
l1U42dF2P1aBlwR2g7+QFr81y3YEmzVqpFEEch8DfVv9e1gyrUwpThG2FPjhYBKFVjcY5tdT8Zqc
7tcxBNcGdiULQEkcLaUk6xTvegyVgpOmR+Zh7twaRmhe+Sa2BUCyQQnV8JsAFYgXHa+1lCgPnD+Y
q3wSWsL2z72+PbMrbJ58zv1HV7LCvpMuvbA+uIciml+UStp+u9Txifu0Ds5HU46v66WyK4Pm2Lhf
9p3MlRWVVFJzHzjylA7aXLjoO+hq9LhlZRHP00dlQGkI3QhMKNS2xYW/A43d95RivDLV638WKGZq
6UZokHSvdTh0e2REy1unJkxy7Wr0O76PmLo0C7Mb2A2OiyYtA09wUfvT6tcLooLK1sq88b37yeek
tJNNAvGFSM+Q3AVYQBzA1ywXyf8ta4T0zgvKQuZOO+stHbphvJ+P5Hgs/wwkBBUlnXlZeh9ncojM
hEWyvn9qkRJR0g/7NuN5zKb8+LsIiEOoI/A28uCba7jBSnQ5AoqYQbXnH3e+TqFTT2IwyYKns1wx
WLDahQxt7GdJgApImmG9jZqukfYsFITHTNBIHUn8p7UXzW7QM5GJrl2kYrMIntGyB8bxQzSeSKXm
2aYGG+U4KMmrSgtzZ1V7povQ+OATleCzEcKwZA3EvZTn01KFbg2s4POKdXJdsKxbU/lXM7UPbUVo
qW/TUV7Qy7ya5Ez8gS2cJqLX/jhxjGVVTNK7P+5Kh3UalHPbQyuWmRji3004P+hkOFSsf2/qMy0x
Makh9R7NgOZPtTdgcOUQ62lYaUUSee1QHsZc+pWwCQ1OnnaGoJ+SyTb03xaU+GaB+53npaYkE6Lt
hfo018XoohormpZiO2So+SIxFvR0weIqhxnodXmRP7JX8VOP4oL2Dg9atX649ShYELO4ckwz0rWo
gEmMg7n6yA3LMH630D51gCpAw4gEiwUM8whNTc89sxUVUfLQyMWz87EJdteNKF8G2CTsNUrxOpdW
miJgYlCheR3MUyTuzpkHgysTKZOhspPBw/ztR2XMIDexW07CPc+YjD8Gy7JNq5qz0G3D8mvuJfkQ
wYKCCietONHU7hTiHnc41/fUVIit++Y2vSXNTgjSm5wQpn5WEUx6/0AKcxA3eqR6pqlDMVafbaec
VV5VWudoCTuwkpNiP6TGAodBhUlPukvq7riQhgESLeLtgrvGuFYdot8Ce2rRKP0GAYpV96Nf7yA9
XKhe9OudcHfRGI5CVnwDt/FpeYMz7G0RlPYcgoRd3+8jCPtYzF8vZZ14kvAxHP8pqBveHi4khfOz
RlNClOOGYIcLefutszGf6zC4AAqxXPTrmjpo8jCj580qhK2rEryQGBYvvXeXmDDzuFFe2FzPgh5n
3Pe76KGbl1EW7Ki0Hv6AMv1nYiULAvULRqV8KlV30QZfsviM9Piorq5GF+gcVIVBW5EnCMf9qIO9
b4gOp5ntuCL4dPwpC1WWPLO4k7va2Ihb4HSmrg/KlCBBJ8a9HkergtGxqxctCYlXk0Z15JdhAZmk
p6JoUusw1H3xfxthutNEf+sGcIigx1BFcj5D+Usjq46Y0eSDvH3uUulwKAtuxLdl32sjrIb5/VMw
T5WvIGuSMiybo6pYI8sJdwI00BRPxjLvrYeZ7kK4p/zEBwegdRF6EqizAdk8qT0DBfZySqhD7S33
gJubaJXrBLhvouzbznF7j7/JnOme9bsOxaqrecY1RQOb7dGFfuVkPUxiOlOnIrU+YtIyp88qIWy3
9VNyaTvjoB2T3CxPM80NfCGxMLlr6dKROuMzbz7vvgJDpBorTJ+iZlg8MYzBFp3IVRH5rpChtgoy
iDutWhuab6/8Z4wqOeuK/VBhWpVdNq5urvBceNmSOjrn6H9Ze2qPIShqW+22PQx7W8JPC3picr1/
XNJl8Y4nO6SEbrqW3fIm+uH5qqLzZMn6AW2SorQg9YQLdevszRMD7xSoOMPwegPMGbMo9OBREnDg
/6+8+XVodct8q+ITJj+eyXwDNLclTlQIFh+DoEqqQ+wXROi+fmfwp+P+jS71ZvuJ2dZcjv3dKtBK
JzQRvAQAuoMJjlyxqwJgUXGWH528iZB+cDNdCBQolFkYepZZ1+LEW0ln6BOKaMr9K6hpusM7H4Pk
2y/wKLKp519tq8v0C5MbES9tOIk3Vs2AbEOrrcF7fjdrb8Nsg++muOSf3tbohOrT9az+ttpq3Boj
t4vh8TgvnpJ5APZIk1hRIvEt5QLthj/k7rXvCj58dQEaGVHWR7fnNA/fKM/koU9HWpFiMFAmAiBh
go2v1Br7bF9x9XzAXvKtT5zWrtuHlqCupOzRaCJwPW+UWh2+CNlp1h3ZptTVicYFXdONovAZfHi1
i7pstoORnJkYhCcXDpuLWcrT5+6cjKzrO24ydBoEquBcqZdeGQD0dlP1lwqGAFJQK0HihNBvX4hi
LL/6KpeP4gbfqECYB3Hc4U/yb3wmEk4huHEJ3JR7VR7Q9rDxIhOudLQn+ejnuH5J+eiKXJWKNsJy
9rVHqgaysUsrtehwY9kNQy99EnVyPxTMaRmWwd+bjSC6oT2LK4RAYseYDNV5Y3QCMpmrRlQADPl7
I+0fIBEZ/WHPQ4S4FP7E1NrwrzLnPeENznsAJeEARYDve8aIrPww3i447CUv2TjyQYoleMqOz3sw
OKiwxrHYgQ03ekoEQdqbv3j81tii+fD3j13yWrqv/ayuRbzPbmXDVdSq1DMVzTmko23k+2Lort9L
pDLd4RbUnoXj15MxjuQxJnYXCq1XOxf4pNGsYM/Qi4B5et5Lpn1mZuqhAw6uABES0uL0t9/5OaD1
Jopg8+PqSalzHpEhO21+gJJtBcarR239LkhP8qfITgMW5McLv64xch7vhQ1kAxPwpys6bTGnAMs1
RzG1mAlxLdeoa0kyVfYqPcyUHgCeYEjY3rxzYQR20U338xfuJNpQQ8eO/BeUVxOaWfQZdlz7JOZ9
vcPfoPrGScrnV3oZ7G0Ht6IIblLlQV80/G4+MAN5OChIsK14iekn4CGoI1SIVhaMMjnzupWS5fU0
gG5Vib39bo+cPTuiABUrdUJntAlDHyhjPCb8+WNSsQNtP2RwkrHUP/i5DgXK+Miuzyf+/lGhXHUl
gan72pao1MK2vSTMfiLwJSRCyRIupRKPBGrNXYmY/Fg6oVFzE+3scNzGsQcF2p+Rk43MrxvQfPst
HEPGe8Z89KsLpCsH4gUzIxwNxYSqrpOJQCoFImEoIv0KiEqlrRBUsac2g5/UTvGTGFBOihArTGMe
HprBBNV7miFxUjYV76pAqmRgsyCCXiyQDOktEcHCiiP+D0ZFhBXJuxKrVGYlnqv47wEPGhew33QE
HCXCLvBtag0NThYdaJFxDPPLT8DgiDIukIEuXEM7FLsXzD4uLbCur31UNEKbbpAbh3EiNHMbqGCG
7oG9+jnLcjSaxPTdfUEfFP4lH7fLKnJo7HnnsHwu3l9XjG6KcMxDUsQFAO7n8xrO5rPAlmboP8dG
XTNvbkpfQDabmveqQVM7H9/Cw5vwpuLbpS/FhO3m0rpmoWnWaAzeq3UDDsu93oQXW2Bw7Vzi/wgG
x+XTsKtRM0ERchNRYm44ET7fISi1OhK3ukm4tKlNbHMHPHqYVigAA7nwlHlbupbD+jju2ZR8Hql+
b24LNjmNspn3FppUsUs792LBwS7PTc9H9XOPjcBs2GI30B2YaBSMiF46iYEttWNb8cf56kMovIZO
OqS4Yypj7SlaIhuwRtcttHVRVk10MsmbkuWwLvnFYsVyitUKXkGcuilwbuOITuyEOCeCAVDZSSuE
ShAWsaPJyvMpeVZVnitEPtILp9ESrSVBgEAGJdnL3mPPHJMZljKmGY0G5NWdOMK0+G77uJICpGHb
EuS/OCipaJOh0hk9uWjkKDlBjqzz2UeoPA47ti4BFflUet2b0qoX8Fe83rencX5BVYki7avU26yx
w6UvSq6dgTeSGlzdQx5DNgIn6OJpsoP3RQEt8g+pZ6cGmrR2R3DTxkmZXexlHmtuWTk49MrUETnR
ymm56ciNr/ei4SswU14r9AAHWLeiOyINMTmpVYUXuzV6Q+o60R7kKz0oeoaV8rPdOp9wI0k0jBy1
foqr4w2mnhqivOc4u0rlQ45x6TOzZozXtU6IUzN6/U7eGswezyn37HRjwVIHzE6+ArcPZ3MCWIKG
ys7z65dgSfkelui0LUN+g85EK6Ar3ROLC/iajMduqz6YdMY6R81+t0g3vAdvOlFAnM/YFXZCYxGg
uoF70SHuWnq/7o34+LIfzwe4o72bGepLJwqRSA4TRD6Iq4IzaYSHIfTV+36MVGh91hRd8JOhyD2l
nE1AAvg1HNRdNfuGXCSULbXeZgNBfMXXD5FeASKuGi9s6DJUhyl7RdQE+zW8IwN8Wbv77YJZj9xU
IB/11RMd3Vts6YrDpLWKxrampVlVzlh/gIXZ0p8Yc2ea0dgemTNJx4qxRZplJYQAcAbgPD0uWzSc
0FRQwyNlVJEHElIrN2BbE3ZdpcM+ffAGURbyLZxuNnMvmHeiHa7Eb1wx6PNQVoSvDI4BIG+5xP45
g0gIf1tu3Vvwf1PZVI/UrrqFxpIh3fOjfSOv1zj+Yguo2UDEsbd0YjfVETtsun7uNYe2I5mtTcmQ
YxazEP5+tP/55a3gE/rOKZyuisVaY+SphVrKyYP37Z5Piuy2180OnZz6xzt84FZsBK1izu215X2i
y+6QqFFWoViuMJnPova1ZHt1XIQH34KRm5+gYqIybvESkpUDWaJLBZ1DGQdzo5xnc8HZ3Zx1Y3wZ
F+7hFoakT7IBKZX00PQjNUXZwCMJbsNIkkYrwy9OhuClmQrwoA5uO8VrohUa1vlpclqmZLiUQMDS
VeiAI2YqZ/QSTTRl+cL1NMXNxLMH0aMueZEnsNoHKOjfKGCr74coetWr5kaHBug33DkfRzneSoi0
nJcRaZlI9/xTz02omAOGaY0kKDm347JV8R9SY0vnUmWwpmc8q6sBEY+NN9/6rGUw/iIn365VGfJY
+fvjsj/TLn0BammAI+Y9Vq3HtGR962/OXk26FVpNrPJIT3mrZvMKHwZ0Z7XH5adEwptO4qiArKJ7
cBhKAWtaNQ33fQ0KurGkAQjn5b4K0+buFxH0W/ODW9HFYop65pTshLa7PWWZv6ZP6Wawm0TGvhhj
bMfNIAr9ttKE4b5cW52467cu7sqY83CZjj72pAEXznGzhi6n13diNiqUgKNQq017RY1vLxSpBwHw
ycF3FOLuhyrE4nd8xLGSWgt29nBzYgckr/199kp60wVUKxblkaGOo27oTp3QJSwY/uUCj6AvOs5e
K4JjYyJuCdYh/OhPmjTD4FJXLOgVOEoRnasaJfC9+Eha1/44g2SBH2AyPF+YscnQa/pbvsFb4MvA
BL+BmK6mmmJ/4tbV0sFNBjTUhcGd24/jiDGlsI8hDze6fjrqiqSUt70ARVOHG5wlVl2O+MhjHIfg
FTDLTpyz7fryoqwG3EPyk9R1SpVTLR7FEP03XHpSX6dTC3bbcqqK6dvfYC3I8ZVdaJkQ7mZ4XBr+
ZQpQ6VrhrAYBXNtP5xjzduIhH74TZn+ka9rYAhnjxcLbCZdhOLQtfEnF7XkPWfJV5rD6q5MX02Cy
AwSL6sYvj44cBRlMqPPB98nbzoQq8xIBk26Cpk6yGuzVmr+LYUBqGS7PrizBSsGdUT1IZWknE1W4
W7/BRvDc+YR1b5fu1zzhpuEZ9ye5x399x+P9vqquI7RTIJCvDXF9f6R0iIGRENQuVBmsnYh8y+jY
sGMFpR0ST8GwBmnGpJ5LPE4zekO8hLoG5tMgsJi2mNbJphqoj51gplMBunHVylY5U6TQZ7Jdih+w
wPfBSIQm1Yyz9XrTRrcV1V1y1IdosvJFMQKJtcttge3LWPDuPJiPuHRrWypkPcIEVStb3eWRA/Fn
fHHEcQyr9JIZcYBbCe3hjuW9FBkk1ewec/QQVak2W1KgNiP5U8L29cHuluwSJv0MY9zYxdGImvFM
+3GzZ2GOfRuv7+05e0/LOlG0syqIsRty6avomYvGcMnlHfOoQfCxneHZgs1FgNQctMSVQO6+Oh0g
413XIEyYyc2/EXhHbB3C7Q9NVC9y+XqBR+MhBFEVkW/zZb838hl2RUzSMY/quNBJr5rubhyq+4Lo
zKIxQXwYqQa7Jf1/zYrKr4t7cwZtfrw6EPOEqVB/c7Y024yMj5dcTWMNL8CS7a++gXztxMf+BZXH
ndpnGLRjnEiKrW/zR+z9Vb3AIX8cfxLW5sikcublF4yXtKWe3ZPfG2YIlxRjL7J8tVbHVrFqR6R5
xAQu0o+YPRxC8loa1TfFlfxD0DfCsQBPAXHj4pNNl5Rx3XILNxfbJwa1DDD2LEG4ov7Vx2ztPUvh
jEXRk/jHNuQlUtg0/l9cmSG2QzNY1WfYD1cQ6fySa8IJ0+g6KS1Nd4cQNk9Zj+ya0n2Co6Q+/SRC
uaul6QsKohKNm7C2BV7Y66atBIomOSEHqqRqx6q7MqjiFn83HI8u85XvAwpU6k/mLKO0GbQ2Za1y
41EyX0f6Ne5w3u8pwG9ovU4QXm3vk1ejyz3XQvlcku8w0Z4A8qYZLjRGXpLj7Cryr/wWcVVAfoP2
HSgkoOEvyWelkjzBYdN33cmsJn/WGBr9rJfgkaUYXqPXL+YmTEU4VnRX37yXqXwx40uMpMgwMs91
vBrbwAVBe8QQv4gQp6KR2jullbMEpchAs0Qv2yaWfQZb9mQynHKkvrJOyL91gA61qlHMACsXgS7t
c940x2zdXr5FO6NLkN0Dk70UFqArBLOYXuTDGew2TxxE90sotXGdmmpQazowFuK0JrSTEZu8dVbv
aHrEw20zHovjxcS567rw/X+BN4ay1uWHULQoC2a3QFMqWk5eKqoRQ973GxmOFyRrsxcD6VZWyAU4
+qMFX+BqNF/kgqyXxvlgDT0YBVsxBZdgitInvTpQuMnjWR5H9DS3Tdx/09/wLB2AyTWWhRYVxlsq
wZLusLz+KFVx0dZ2LO/3lWoWgSa3zdBtup67yz6c8hwC7Z/0zFPsWvjE86UWsm4EXiYQvJtCpWpF
xZEtA0idK/1z/g/4YYR/+AUbvJthfGFPV8m6eNVZ74RWfZAkbHvu2JZ+Tjx6riQGklthEmrNjHiZ
j1kwgQ1ZqnITsKnKkT2QnPiUS7fNJrMzWz327V3NVfHlELO+ZOuchMKHcuZl5Fa9x0o+4TiCPSL4
NWoI72gMpt327FpPIomToPS+4MnGQk5ZUWTDro7WT8JAsXcqid2Gv9edXOHEfqbQ8twxwLUU9b8Z
/YFgFWXlCmMI77yWTTYWPZzBtTY3awG8+cIJlNTcJZqOP/W6T23lDUUGWNB2C1ykPcLLD8ZX6+1t
HGyaln8RjOE66i/SReSWgKoyYmtIoIlHHpk7CUYuHonlZqNDYbjaf8jVcuUZ4/lYe2+RUzf9DDaW
0a4KKJO5ORXPVsVy2vz+QztyF5mi5zlBgzGysYVXjvMVUQ5PU9CvwttnOqinAmzItAgEGydhHGAf
jxcWs90bzAwGdH8/L74iAyr4JevrREGjLCTpcOg7GBiO5l7lSZlkqaCWY6o23L47TkV0k1bSZtsN
SLkLjWX3xrtBsaPHdKty+JY8yCGbTR0H5Y7DNPqDhKm7IJCqewlKLodDdXQ6TKCi6BfrEFrzDarU
hVzeQmPfFtzRsbW0lkjqoh2lhCR+axoO3+tTFA05sHE+RitTR3L8q38lUh/w//znnPNOtpPOKzCS
K+EWHNo1EluEMIFqod/6vLtI6GcGkDxm2GBYzceuxqMawHTBwU3Sp9yiKa+moeA08nSTN+otjb6O
YSTIGm8an4bWiTlidNc6SrNjX1ceQ0I7juiSYSMI8fbGv0OBrA6xuW+WKNh1xhZUvWXghUfj+o8N
803SsVBzp2mMLt8yFGUt5hzc71qb97by9n5XhcN3+2LtoF9ABWXRK57bHaF5d3nHUTfm43Alq/77
UKh6/b9xlZwFE1NV9uNYEebAqfhr71+gQlWbgWjyimHvVJgTbFe9u7/twDGjNv5V+r8CqAbE2pBw
YxFsoxmU1gDAVXxISANWdfisTiVosDkyocruiOtWzSlIi04Gs1c7XdvfHYKldMk5goKks8oF1R6U
CbkXKPluurk/sXVcO/2F2Mre0d4K6WpNi/tyFLARjeDhPez5qBN1G+9m/QuiN2cPmPKeuhiHuhUo
/CNQIfqPwiPcBhgPo+G3gp5e/uG9YRUqdY+XTrr+rJqCvSUTuv1aqZoo3GEz/BbhUe3u4AFId+r9
Z1YdLyGQKwuycPjgAhQz06osw/UnbzOEysHFbNSpjaMgfWUjW6wFSW+rGbMGQzbl8Aca6qUQNZSg
DIRNLYM53UjK7o8zr5PwKMlDUHynbo2pvtbnjBD/3lcg3WuFy0sM3s4rntcaIAncYMdoWl4Wb1o3
6SUCtfqBYqpC3mueqz8eJvXXSInfMjHouGj4Ne6lIxPrAwva1cCZ5Dszy4bOl1+nokWb+gqp
`protect end_protected
